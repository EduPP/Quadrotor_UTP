  --Example instantiation for system 'NiosII'
  NiosII_inst : NiosII
    port map(
      dclk_from_the_epcs_flash_controller => dclk_from_the_epcs_flash_controller,
      locked_from_the_pll => locked_from_the_pll,
      out_port_from_the_PWM_1 => out_port_from_the_PWM_1,
      out_port_from_the_PWM_2 => out_port_from_the_PWM_2,
      out_port_from_the_PWM_3 => out_port_from_the_PWM_3,
      out_port_from_the_PWM_4 => out_port_from_the_PWM_4,
      out_port_from_the_data_tx => out_port_from_the_data_tx,
      out_port_from_the_out_test => out_port_from_the_out_test,
      phasedone_from_the_pll => phasedone_from_the_pll,
      sce_from_the_epcs_flash_controller => sce_from_the_epcs_flash_controller,
      sdo_from_the_epcs_flash_controller => sdo_from_the_epcs_flash_controller,
      sdram_clk => sdram_clk,
      sys_clk => sys_clk,
      txd_from_the_uart_gps => txd_from_the_uart_gps,
      txd_from_the_uart_xbee => txd_from_the_uart_xbee,
      zs_addr_from_the_sdram => zs_addr_from_the_sdram,
      zs_ba_from_the_sdram => zs_ba_from_the_sdram,
      zs_cas_n_from_the_sdram => zs_cas_n_from_the_sdram,
      zs_cke_from_the_sdram => zs_cke_from_the_sdram,
      zs_cs_n_from_the_sdram => zs_cs_n_from_the_sdram,
      zs_dq_to_and_from_the_sdram => zs_dq_to_and_from_the_sdram,
      zs_dqm_from_the_sdram => zs_dqm_from_the_sdram,
      zs_ras_n_from_the_sdram => zs_ras_n_from_the_sdram,
      zs_we_n_from_the_sdram => zs_we_n_from_the_sdram,
      areset_to_the_pll => areset_to_the_pll,
      clk_50 => clk_50,
      data0_to_the_epcs_flash_controller => data0_to_the_epcs_flash_controller,
      in_port_to_the_duty_1 => in_port_to_the_duty_1,
      in_port_to_the_duty_2 => in_port_to_the_duty_2,
      in_port_to_the_duty_3 => in_port_to_the_duty_3,
      in_port_to_the_duty_4 => in_port_to_the_duty_4,
      in_port_to_the_entrada_ac_eje_X => in_port_to_the_entrada_ac_eje_X,
      in_port_to_the_entrada_ac_eje_Y => in_port_to_the_entrada_ac_eje_Y,
      in_port_to_the_entrada_ac_eje_Z => in_port_to_the_entrada_ac_eje_Z,
      in_port_to_the_entrada_gy_eje_X => in_port_to_the_entrada_gy_eje_X,
      in_port_to_the_entrada_gy_eje_Y => in_port_to_the_entrada_gy_eje_Y,
      in_port_to_the_entrada_gy_eje_Z => in_port_to_the_entrada_gy_eje_Z,
      in_port_to_the_entrada_ma_eje_X => in_port_to_the_entrada_ma_eje_X,
      in_port_to_the_entrada_ma_eje_Y => in_port_to_the_entrada_ma_eje_Y,
      in_port_to_the_entrada_ma_eje_Z => in_port_to_the_entrada_ma_eje_Z,
      in_port_to_the_entrada_temp => in_port_to_the_entrada_temp,
      reset_n => reset_n,
      rxd_to_the_uart_gps => rxd_to_the_uart_gps,
      rxd_to_the_uart_xbee => rxd_to_the_uart_xbee
    );


