��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F��J>�����>�����HU�k;�� �[�+?�w)݁)��>7Ý�4�B#�"u�%��R9�*2�	φ�v&�f�UxJ�%�����OOL�mF4O0��%�O6?][��W5Ff�i�]�E҅u#��Vg�n�����g9�#���>rh�W&��zCu�M��{����,l6�`I��3����
X�	�@�#��꘲t�}p�ũ�g���.�pæ�dbB�:�`�(8����Q���E�m5���[\[��Z�Xe���z��e�ّ̀�4��'͐??�r���4U��e|{��s�_
���^��5���ЉS�u^R��r	
 K�Ԓ#tO���?�M�ΟuD�(}�G���|E�,n���;��"�z���+�rW�t�ǟ��[�z���Q��Ƈ�b]e}s�;�H�:��(�=����ݺ�����)%����j�⽾I���G6
�<=h��/�[m�S�\I�.4�A�1��S�S��h$��Mj�1�~�P|ul�P�,hM����R2��U�&tˀ.?���9i|������u��F_8�����-�'zx8�~�$	�	+��D\ߍ�b�+/n�f i��O>U�9���mx�������V�K�`?2_�ĥ�3?@A�ʺ*��P �j�C�
����ï��b�A����[���GE��\
���k:
�@�fv6�xR��G��� +�U�.?�T�:y4�_,��7�&��!J�+9?[X��b�1�#���l��;�l���@�7��-�c�)��(�E��V|��i�P/��0��9���E��bQgb
�fYR�E���Do5�����6�r��"�Ҝ��9�=�N���5�Wؒ4��P�bЊ&x�`
'�97^�(9�!W���Dxp@p-/��0Iﴓ8�Y���v-qk��;�Ң7ժ��ٲ?������TH�A���o~��pI��<C�@}|ل1�ў%hz�&��-p�n5�,I�)3�����*�}{�.�O� qI�naG���"0Bσƥ�pl?[� ���,.χcFP��&�?uP��
����������K�,��hXJ��Q��^�M����ϕ��< �����d1�r�UK��c$�;�*�����l��.s��G��G��9��H�Fdy ��M*p����|��T`��GZ��{��4[�@��v��yq���p+ے�5�4 �:�/8~/���E{ЄѲ�1���F<�=w���$�ܛ��;� +�z�SqS���~)�g81m8{3�!���rJa��;a!�j��h�"v�A"�_+S<��'9S,���)��G�x��?�A�e=���}��#�7e�x����vj�)��'t�/�d*��J���[k`��Ƽ�Wm���a�Zc�u�A��a�jM?���b��d�*�['����Z/������mEӝ�b�u�"�,
\�2&�g�+�#>�B���+��5�l����/����	@Z�A��r[�{���;�U����y��8�zY���_k�M\+�{��TÏ�Nd���H/6^�~ub���}����M�K&]���r�ͳ�� � ���+΁�h���v�bU�� �����!jE1��?����J2��Al����5��#�y�ؑ��'?�B�M#���l~��#h?%�K����D���*���6��/t�ɑ�s����)�i�Pv��,H���]|��-��-��Gxsd;D��V]�>�5EE&)�-c��9��7��З�`	_IU鐎:I�F�&{�,CcdU���Ґ=�g�p�uus$�O7�/wL��dވ�{g��ei���҅#��p��B�&��d��%���Y}��^穁�2�BW�C�������Z���yČeM~���|�Ey@F��4~﯋2RY_*rb���0S���
6����Y)�&q�`��ώ�Y�7f<�r��k�f8�%�Q&_r���.��r���;o3E`�kp7��{��G��qdIP*4~�9�W|���	o��4R�����(�-�-8K�������Jc�G�&��B�>�N*�����2QP@o�~�ܬ*��󬏷��nS�+oA��9��%�p�A@��]��h+l�?9_'x�5��g�E��"Y9�W��C ��(Nb��Q$�a(�d�O�Tͭk�ꔣ��w��;�zZu��R� d�wf&��4�T2���L� ��w-/C�喝��l�놞��3��L"ś.�Xnǖ����_�;��;�����/	�O�0S�/w�Α�&�b�y����u��I�U��2\������U�{K!�cN�0���YX;8^&6PD�ߴȓ�b���~�T{�ْ2��]�-� �^f����B���?����JFO�O�P��c.|�!},d��W^�`�:���ȓ�U�͐
��ۥ\�+�� �����ݣ=���ӈ�0�)r'a���s� Q���eTcu���4��[s� �C"�v� ��p�{^u���4~�us�1�~��|����b�����s&������@&���'�)u���!�T�����,ћ��Z�5B_��INh��uB%�q7�_=�)H�3�� S�Єo�i96��閳+��f�
U�U#�v�m��9��6q�y�P����|��]U���h����@��[Z�&t=�'~��������!rB�/*@��O��	M�qf�.�Ǖb�:ge�P�~B�*�8�SV'&J�t�P�'��M>��PW\�a��#�g>��HyAqHr���R�d���P��������.��nPu��޷�=|?|�U�
�Өp�T����zMI�T)�#���rw��4��X#�k�tI$�ʼ�%݀@|qi����l��iT9��|[��s��h:�����+ĳ� >Ε���N������8�	 �ݣ��oԉ�Fv��M�=?ʥ�"��мb�ZT��zZ��Z%��jl�4�� �x�5�1+�>;�{,���Z� )��gO)ݤU4����Z(6��D��^����l���`U.���6����L*w�P� B��R���%G����z��Ϝ[]�n1:f����,���|F͂�p(Zl�G&����p P)`�yG��C�f�=6�=�A��e�M�(/x|k���/7D-ŦGY9`�o��a����� �K�d ��7�8&d{��D>4���޹B2<i������]��l�-��Ӿ�/+|��m���+_�.͓x�v�;5i*\1͟���E)�X2\'�����{��߈�%n�A�����(u��Y��M��(&�+8�їc�K��Nk`��Z�5b�F�UD��k��7��g�-��㋻ΰ�t��&	��P����%��� ��7|"����Ri<(�`D��p(�:a�+g�����lW=�D������/��zyw���SV��VI���"�"������C�Vf��oҽ�,��"��Z
�zq�=pW���_��c�F��#��}�sTo4���(��٥ ��k<������������GO����#�I"^����v��
#�N���7��9������X�>FH$����U��u�'y(-�d�?w&/>7$6YO?�U��6Y_(�S;XC����Y����U*]ڃ��b%rJ��7�s���Q�|%������y#�*�;a��$��4�a���*쫺����~��ix�i�F,��5�k9�E]n���&�.���|m{�m�Jj�Q�� M��rm�W�O�Nۜ�?��u��xY-�N#&z�s�B�)�F8��^^��BO��ҹ���#�оԒc<�U��9y��'�@\��[K�F|��@��QI��is3mB�n�f�wmK���YA��VV��{�l�أ���p�=k8��s���ecޢqb�$���)6���ɼ����{�Ԋ\������Gn�G�$�VZt3i	��oˀU��iGP"�=����J� �=���H.U#��<�[������X�y�I�<��I��כY]�|۷���ɄJ�H�q� A�R@��nrO����>��Ϥ���L�Ue��g|!K�q�߯����[p�c�+���/�(e��5�ՠM�,`��F�@g�!/���C��oH*x|�0�?�@���	vz���=YN�B���~�� B��/:����f�_��cU�J��.޺Ō�+D�;���=���v�+3�>ĕ7/S��ݒ�-��'a\��R'qK�I_�*V-���56e��׆���<��{���e�&1��e|Te�c!�B'.[�8Bq8�#��$�)3�))*�'*'o�U�Tb�
����.o�I�g�hdY��R*��h������f���^�O�=��E���0m�`�H�wjt�[�.U?���<��<�u�u��F��NO5[K���O�g�����G���(1e�d��x���=�#�v�D: Tc�5��y�3�_f⑂<dK�.���N~�Z����Ð}G��m��9�O`���阮���P���⡳��=d�����?W�J�`�_oJ!39��2�8��@�������z�YP$+�Z?�k��j�#}(�.`�a"�N�g��k,���N�����#�QA�7�x���a�sf�c�k�g�����S�8�nQ	��dA}�_���g��qH���}]�g�+�"��[0���8}�2�i�:$g�����#������?J�x��2���)̥,�x����&HK�d���n�.G�G�3�~	�wv3&���Χ�6�?�Nlf����!G6p5^hr�fW��ׇ�I6c�� �0��`��q�@��u��MR���Ώ'�[�$�+�B`���*,W~^�X��hG ׽����L����I*���C!ox��m�����D�Esr�E�;g��N�!X�[��ߧ���-�G����`T�A�"W\K�B`P~A|4 C�r�2Z7?�"å$�J��J[�=�*����՛h��p��m�j���GD�
K����j�N�"Ic������C��tf��Mi�2]~p2�#-�Ҹ��Ɨ�r��ܭ�v5�q�&�ށ�`^��	�X�ͧt'����|��Z��|,�i6��Q�&��4Yl�ڸ5a���f��Cèik/�0�,^�:�ٰ3;y�k��,
hq�9����;g�N�G!X�*���c�M�<4�0~0�����Џ�bPN��6H0:1�iҬpR�r5�'ǘƣk�do�*Пܽ�N��w�u|��x�G�v*���܂W��%�����i�h�s��Jf�C��ob����*a��L4���^15�!/��9���e�p��/��� ����]��:��.�D��6�d��t~u�so���!��_
9G�~��qt����wc���uM�� ��\͏�M1�5Q^Rˑp*���$�~��R���/l��
_.����dʿ��k6Ξ1v�5Q��������?{��}�:�]��*"�kS���b������;����!Q�^�	�������>0!7{L �uw�[�G����������	�/;�6�[��)��M�'^rXs��%�IF��!���n\ؖ�h�xܡ���e�h�p;���@��[�;C\����Y�-#����Dh��p�IƝ�d���� fl�?F��M4���OU�����Yг2;���M�س�����Q�2�2���E��x.�1��EûJb��<O�|f#+��&�����\v�g�7��?�����K*Q��f��и����	&��w/�!p}�>����Gy��	�K[�)���j�ݒ�\�gٳ�,����`��a��Gҁ���zA�`���2)3�f�$�P}7��� ��g/m��'���>��H랢m�]��J%�3�V�3>�r��u�k���A�����i��)R]t+u��#Y���L.��0��r�&�?�j6P@�`���|�8�v8kj���yc�1�v軱�}�LŚT�^�f����;PG&گ��a���s&�.���<Ie܀x���;�� i��ptUؗ��6��P��5'J�2����R��uFv ]�uޕ�H r��!�3=�R�e9O�`�5�)Ɇx�e]<�{���kc�\��}֒���	9V�j�ڃX�C��9��_7lr2Ql�Q�6�=��Dg�V��|=��PO0fct�S!�>j$��/�M}��K�ef1(���W����^��æs/��t����&s:z����g��w����!ɝ���N�L�WrK�&�o��W |�+���S0g�)��Y�Ɣ:/`n�Z���(�l���3e,��S����x�6��X�͍�Ș�*���JݬR�8���VZ��2k���
�A�V����T��)a�fGq��Vh�r�neM>��q��(�o)b��{����`cnR+K9)�t+��K�o�����d^��	�}�䌆�V�2P�`[�ʍvn@/�:Xz�ڐ��\�7c8�n �{,�ql5�������$`�ȭ:����7��O+Ge<������(��Yո�n@�`�>s����S{�j�	��r�@��F��� Q?2'4iZX�D��M'�C�[�ya��J&�����l��Iܧ�Kcݶ�TC6��Mn
�Q�ԗ/7ǅro���xG��-ȁ�9=�*�cYY�w�bc��a�j�[N�g����\��k'e��c0vf���e9�b�K{�M��m�EGńƲ����
�W���?��r�	��_	� �i�$<�`o�pu�� �ˍMlL�z.�=٣�QL�L�t���q=6�JO����7�B�[u}�ݨ�[=,�2�ѧ��S����!�J�ެ�d���/��!�ף�4� F9~�����m�����X�m�ydD����j����{0��s��\r�k'�zf�9lS�M�-Ά����|���`]n~_/�8H�g,��F;S�Vb��H�$0p�1�&�o���^�?��4�q���퉿�2R�����U��+2M�lZ�'S�=��j[�4�!A耓B�+�u�?`^�m��]	�xۉ`gwY�DS�3��8 �w���?��eK	\ɞ}qxσ c��:�� ��/�߬e�ի��|߲������T ;>]����X�V�m�6]� u-�}h\� �t���
�Tp��11��4t3���*ĩb�/�Ż>K
�1N|���+�/U�%�"���jո��G��A��vI���@:&���2���]��w���W�d��5@dB��D0�9�,�O��6)z�H��T�w?j2�5�諙�v�n�����ˈ� ��-�JS欣�|�HU�������姌ՓI~�Ft U�[5���0����⠶6e~䉿h|�8� Vl��D��W������[�s���X�%P,t���\�f:����֊
}p���T%뿄��a�9F��sp�ܽ����yנ6X���ޑޡL�edoSRZ��gR۸&k�k�������~^�[��L
O����&�ڡ�%��J�i�d�ͅ[ѩG��E����0�/Q��e�h��A��p�ҏ�mgTjr��o���$[������C�FL�1"D�\#�b��6ƞ���d��]�v �q��SG�~�p��7�,�i����'vK���M:�z��C��Υ���nZy�h�s�B�����8�"����`H1��ǳg.��߲��r�瘪'�"��,���z�Y�~Nk/
��vs
�`���:��ԗ�^�q$�*XhKD�Т�a���N��L�?����=Q��<��p�\����1U&l:܈�^���^A�ˢNy3I 	gNߋ���M����l*����c�3�EnQP9������/=�^��.T˵���S_;��y���Q+G�Z���/��ۧ�Y��@$�|9]eˢ��#M ፱}�ZE��Y�Zs�L�����Rp1�V%ʲ��ۓz��О`Y��܏��뫜ɺ'2��?^�զ���)���7znJ{ض��nY�.�D�?����ǝ[�}Y���Չ������z/�F��c1��I/h�S���X�b����	��,Nfk܂�%��(	���vι������\�w�6d��Ϝ��Or�ۋv?�!%�4��RhQ^�[���\P1�\����K��4�َڟ��t�C��ݓ�כ��18�ΕG�9E�G��;v&�����6ƛ����:"LK�"���,�����Y���u���Iә����0 �����}N̖	\uQ�X��sZ�;ŀ5ٵ���*W��1N����� UA4�Z�26r��S�̗3�R�y��Ժ<�g�^�qu���:��:��z�$m��
�@������=t�+15����hd�iখ�4*p�粠}|?�FS�Q����8��(,��L�� Ȑ�^v�'@�<V:»�G�Rw��Ւ���������o!hK�򸡞��a�o���D�!�;K�+ٗ&���"QX���bZ��� Db�������^�n���p��?�V]��J0-~]@)a�F�Ȗ�JIU�pT��P�5��O����g���7��ꈎwS�N��8�Dnpc�?Ǌs�`�k9�z��"�T�t��a9Y=wi6����M��x�bn;��hX:H��;_e���EUCEz�m�J����՝��������b���T']!*���Qn���R��R_������$u����,�E���X�?~��R�����&��K(OO��A.�HC(+�@9��:�W@�5�!��gg����P��,����6VT	�ch%��ހ���ha����u��^
=_�- �y�����X�gIW����S�u��=E�8I�L�0�h�S��a��)(5S����he	Ql�xr!/l>�Q���p#�o���������B&�.����%喬,�Z�p���6��B��Uq����X�E���	Y� W�Ɲ���ꗓW�6�ku�z�AI�%�_����f�(�Y�@�j5�2�]kMp��%=���{��9������#ٜ�!�X���ý�ы���0�W3�!]��#<���v{��{@�9�%�\'�ۀ�6;o��^Q&���|�����{W����mS���I�fz��v[�έ�ZT�
�@�O䆤Qvw�6�W(Ǹ���X����R\�a/)�5��;%/�5c
�K��prSF Ut��uL��SVA[y�&1oq��>ēVI����A���׹V�%[I��aMGފ�\�;���ͱM@�x���/�3���z����m?�^���乴����l���	l�+�	3@�BȽ^������%k
�ٕFMW���h2�\#�X�r�:�;�n��W;��^Z�"�)������|���(T�k�㢘�����jWO��-��9C�����7HB> �+���beGo��4G ��D���:T�z��@��~ˏn>�e��3X��3�&sGi��f�������p��@׮}�QP 	c�[Go24��?o?g���U-��Ưk��0�h�׬P�iY�*��tj;/� p�����a#���7�������3���9\����$�m������Dfzr3�ٚ���6�҃�ܯ����S��k�TҒP3�(�L&ܺ��83�w'���j�5����d���e�:�?�&� �o�x3i30�B�ش|L����&O$��Wq���Im�X�~fW��e�4�cs�?�,Anf��%I&2���l��_u@T7_����P��:�^9��ǯh��(�VH�G�~c?V�_3if�HQ��V^�7��ɖ�����{�o���V!�ӵ��b�7��[ 9 �<��G����.�ao�t�fY�&�6�lf�$%��4S	;u GD
�:@{-n!�I�����?��~2zg#�ҁŇo��<��$�t?s��sA�o��c��������� ����U�0��e�C���`w�'�GB{l�x!z������=#
9��o����R���;E����~�'W�O[�0�/}�ˢ�����.��Q9�ubF��%|�ʆ9�4��m\'��d���3���Q�.C�gu�#�Ί�˺�3w��75;:�9�˸[����ܭ0� ��|��趃-X�ɚ=���������v1L���r�[P9�Tr���?�Fc�v�Rr�.�jx�H�(���gj���d��q����ŭn����������x}+ �a�@Ű�Hjb�-��rM�>��_�K��Aܚ��5���N������&eZ����%41�=i�B�
U_�Y��\��mt?d�#��O�%��w^��i�� l�7K�>qFz�/��(f�Vu���K�K)i$|iS(����Kz�
�����k�~�Z~Qs��Ό��r��������MV8��t���y8"���a��P�����j�@����t�C��_A�(S(J�B@ŵ�X/�N�y�{=��Jop��<Ȼ�0~������zMi�{kewcE(O�˚,2y4���H��+Z��n������ω�����6�NP�Q|�����O�MLD'����J qHB�����
� ��1w?����`� �Eg��}�/4ɪ@2�=rׅ���;�)�8���hH�=�ΡO���E@s�EtR�[��Z}-���2�A�}�m:�,YD��@>�t릐�'$L��WS��7�F��N�߯�HN�I�.M����Qu����rht��Et-n���2)���gn�7u�g1ED���6��5M(CC�eЋ�P��~;������; X�"@��������JM�������	n\�A��Ҿލ`�ӝ@�F5��("iV��݀�|���D���;gfҭl���A��� b}[p�M���$��6�zޑ5�>��񗦑̡�u�5h��Lk�BAZ+f
�ܩ�4~�zn�`����dC)���"��L�.�����bl�?�G�������`8%��0��ր y�?�ٝ�銴���N$&��Qͥ:���ޢӷ��Y��CQ��˭S�V����� ~��hD�F� `�h�/{K�/8ߌT�?��۴�7'�l��}l���'<h��cVPb�a~�u]�-
���~�Ȫ���'۴2��UR����N��8�rH s�ש5�Z;����@��؇At�pL끵Lx>c��<ͦ	���ʢQ_�$��w_�s��+�`(�x�]�S�L������1����`7βg^��b�����}K��>�k;���,��m�4Q�+�����Ă+ d��񄐄�Ei�UA3��MB-���4��f�E��d-#�RXF�~���P��kx��e�Y���w̧nS5��������~f�K5WI$R�8�$�7+<��	�A���9� �Դ�"���e���/B�qUv�:�	��rr
طPc�9Dy������7�'��-�|0<�c������ߊ��S� �8�8�|�;Em��:D�Y �0�r�5P�"S��5gN����a��y{�|˞y��SD��ܖ���X�O�'|��#M�^%|�!�����庒*�l�J˖l#daKL%�y�b��񛜖�����P���)�X:��c.���̔�W|#����s�ڼ���m
��/��Ą���j���1�K;aW X({�=��]�Ax�I�Ɩ���$��AT��%l�ѷ��b�wэE`P��0�O�-]�ơo`9���;����%��*�/�����z�C^�U��?o�m�0��V���A��AH�����բ!A|֚�EG�P2 �p��k����ovA��F�e��7�͛�F~��?��#6�p�w9zV?rq;�J���Wk]�-��(
!�|3?���\��5g
_8 �^��*ߦ��1���-p�^,�TZ���ڋL!�#�ˤ��囲�����Y���Ь��Dh6{��C��7��@oT���ѝ?�{���X�w��ٱ׀�cS�r%��?h	xk}��~74�6J�M7@<Ϻ7��2"rA鋔�����8+4i��7���}{A:�5��^W��'MO�z2ybQ���i�{�]YX�H�&�X����&"��8Q� wu-��fGS-�Q�ܒu$�-�Uu�(W����B0��,@����IC,V�'Ӧ4|6
#�?��}y���lF"�]��W�DCV�
iІ8��J.�u�>�c���\u�����ؾ��~��O���0�c4E�kB�ZLow	%�VlO��b���#�>L��c\ q{�&�E�O��ްo�6�&�?O��_<a$��ÝG+��e�5��qK��c���U�p�)�\(��7�5��໋A�YlH�4��>���T �r.ٱ[�$�ID�[��� l������} ��SZ�YY?4_wن�b�J��%6�^�y�HG��S ����L��e�YI#Wu�,�:���n��5l�����G�g�k�Z;٧�|^G�$��W��;m `���^cLz'
����O7/W��'�x��)�=&�A�LCF;�M{#�1r�nͱ��>�\�>FF��h��������e���pU�6�_ʌ/rh4��q�P��A7)Ohm�FEu���|�3ܖ[��E�A/&9{	lm�](�<�o�ܪ{�>~��3��#	]P��"�w��؝���I�h�K/L=��@Eک ��;�+�1J$)���;T�K��{KU������UKF�{Dȿ�i@�Td\�x���7���4��dNo��wsb��}���{�q�l�_L5��	R�(����EJ�j��U
Ә�"�r�\�Ү�_��]��<V���@���g�����s��qL1��Za��;�ƿ؍�#$�7��ȓ�E�����a�Wt��ВE`Aw3.���:��� 9���hl�U�@,CM�,]�� �!J����j�t{��}�=����
�Z�|d8�.�G)=���.$��=;Zvk��TA� ��;�gc�i�E��%t�+>H�,-�����ץ��ޟ&��<{G�c� 6/�ŧzAC$��te�������e�Q�:t�y ��D�_��� P2���l>*��8D�ż�CSQ�g�t�#I��A}�!2Wh5Q}�1���9�ۄ��K>-�z�0�!`|��:��	z�t\6�����Z)3����Q<�!o����G��m�϶��E�ZƋ�������d�_K�Tjƣ=�4
��2(�@���2�t�Gv�BI�E�H������$m��Ȝ�$s�O���Dl�)���x0�x��K�w�mIY
�Y�XC��K@�a�J�iP�u��Ƴ������N�@��j��X�Wz��!�LM/q�/3z��{4(�HԊsv�i�[bsI�/]�A~l�|��6L9��L|x+�e��E�ohp��7�L�9m(F��0?��h�H��r����GJ >����멮����Z�B�]�M���u��,��^'M���"	֓Zُ7$w�`Hn�q��$�c )�w���j/��M��G�̦�S2V�P{�	(?��oUk��� M�W��M�:���A�j\S:�����y��&S�ʺ_�5c�Fϩb{��~@{!��n[�q�/,H���L�j�4��xj.��Ur�A�89\l8�l�Ef�ex���y���A�����t�n{����Y�iq��׋�U(�]�`ڂ���Bﻞ��z��.�������8���O�ǃԆO�a�!�|�l�-���R�E��dI��1P���H�m��ix_�������#�2H��[-�4�;�N��'�;��I�f��Ʒ�O'5��wgmݴ��¥6�*6�8s��^�~����z!�V��N�o��]m�����٢j�.ۗV����+�b�K��U挃8�D~� 0b�	� ���6�/���y'�}�~��!/;�5�����C�
����㵹2R8�2��r<�~��T��-�vn@.�Lʮ��@�a�Ξ-�J�
z!�Ac3W/7�߭Rug�JI�i7&���}%�PН����u`�s@�&�m�ߡ{;�?��w���.7��me���vM�;ϥ��
��p�bxA3�_UZ��$M/"y�Ii}����c�j�e���[K�W�M�����t�A�'1��(��-����Bd7�Ք�)*\5=H���}�ýh� �O��e�כ(��;z��K�-�A��y�6{RwE�/��n_�KL�t�l�������G.�>0�h-{�qZ3s��Y���;���A)/�ug}	@����Hl�ȵ�8j�USz�^2�%���R�������I"�N�qzK(l_��ǒ'}Wv6-��e� �o���v3�p�X�=
U���WH�$u����(�A�GY�3�9?�:��ϡH0QCgo��l�c<�y�0��F�.~&�^��������o���SF��H :o(%�6bG��t¸�9��%��r�62�B�h�v;bW�y�p�exlQ��6�$��)���ho�B_�r�;l�BdO��L���{�G�(?a=g�����g���:r���c �(��0m\'�H�#�"0�`�Ž!��լ��yy�����>���̗��rBFհ���\�IQ ��q��;LLނj>��[�aвF�������f�̭����'���d԰h��4�=�T<7��`oMD]�U�>�U�aw�.��2Hʁ����=4�*�V��RZZ�R�����C�ݪs�%���L8�<$���_���-qϦ$�];��*֟��Hx.�rM���Pm�~)����x?�b(���u.�k����|���A�9�Y����4�g:o"�8(�S�������G?���b�!SZz5Ľb���y�k���ʩ�w�"1W�Y�(]���O�r�\*2����&sf��K��l-a���|����=��`͖�S���[H�[P�M���^��P�Ql��L�p�7-��t�J2,/Lq����R4j�B0Ѩ��`�-�'b<�=�d�����0���S9�A��]$��r!���p�[�V�n���ğ�ET��J���������L��-�	@U�:�,��M��~� �T�C�U�Z�����zD��}��(��+�_�â��c&���k��Wű�|��{c;Ԃ�2�c�L����Ъɓ�7�a���T$���6�=��PH�Jo��_�&��h%�ް;$��!U���^Z#Qs����&��1<�A\���C�K:�c�[�b$3�w�<�'Jg��ja��fK�S��y�o�XC:*�zu4�+��S���dV	�b�B�zhc[/n"o<��C�̮%L�!A��(��f]�_���n^�ؓ����©�
I��G���(G��\������h��F*>��(���P!�P�84�)�3Ê��GL#z�&�j�0�8.�u�v��?z�9�bb�n��j����E�������m���L��gOP[<̣o�~$� ��?�ÇF��LW��M1ec�(��`�VU��*l\ϔm����f)�m7����'rO����>n5R�Z"�d��Pϕ�u^ȻZ�1S������S�$D2 �|������ޅ�=?C�d�Z�-�i[FGr�`>���9v3�����4�u�?e���y�����&_ j`�G�'��
nt����5MA�f��r#���"��a�n���/�ճ�&�z>��Y��.S�Af��=�ǩȌ���Ή��Z�{x�8���{O
��)�C3��*�`�Cϴ�:(��k�_|%a��p��}�V�������/4�h��:�W���	��,��謙Z��,ۣ�Q�O�T���u|х��AI�J��W����~��dX�مm&���9PD`��˝���9�<��T�(9��m�n7�ǰ�x��:��]K���O����}Mm[����̮�$�	��'&9=���"�'�YTgs�v��h'�Y�\.�~
�c��9n�iK����G��x#Yٿ���9֭�ut�zQ���f_�{��[�Xn�44��r�5��96��q��V�&c�M��C}~R �6��٩�GX#Dox�]�p�#~%
mE,��V��d=_�s�����T��=YO�OkI����
�'�&�h𠰣S,�0-Pv
w���8�`<eQ.�P#�y{}M51落! T�<�>P���	T�5?n5<(Zq��->�	��S�s�l��-�,�.�(XC�&�
���Z1�e��U�;���
a�x�_��ޥ�x��5G�����8���ʣ�����)Dl� ���ʜ���E��uR�KV��a��4����VQ���eB�߆�hQ;�}R��@^'�G	�`�������v�k_e�df���s��2q!B�<������g=��w�7�3 8���j��h�.�:}�M7�P'�๐��e���`5�?���qp �1t�W~��u�,�Z8��a��C�+nql<b̛'h��Y� W@ۥe?��04iiIop�4����%�֖^�셟v�Ƶt>ľ��X,y�)�,���f`���B��:5��$��'4�H����n�	�$ [��屿�2��W�m�2L;���4-g��:��n�u qV�xE�2�g�r[k�y���/��T�w��x�b%&MS��s\���=�4���� ���9��u���Bw).o"kxM���`�QKn�[�$��Yhe�W��a�d�R��+!�x���ر����ò�QW�Z�������(�wH���%lI�oM�K1�žb;A�Xx������i�P1Uv9�C\6~Xg���1�	��1��p#'���"�̫S�6?��oin�/FU�� ���	�mI��B���'7�����T� {�l���f��p�[�^��9>s��+ლ�eZ�*mJ�.��Y�gs�����'��N�����r���C�D_�F;�O���j�`�'�Ƞ��9�<�e�Y�`��`�9F-T<��Ad��AR��5�cc4�T.
Ɲ����}�g�
�z�@,(��#m@���X�UŠSe�aǴ�8�t�A^��4&)�� �����Qz�d?7S�g�RFw\v't�G��j�����\3$Ȕd�ʏ�MjG:�T�8RhmTY�������4Љ O��6{���W%�3�ط)v�$C��J�M-Vm �Vp��ڞ���W��_�r��	��}��R5W̵*��ɺ7��k���ip�_7�t�����h��JF����ٯ��qYp�'[
�uB�͜��y,���`OX���<�0x�j;e���ڐ`\)J��Z����$o�W}�+��v.+j��.~��˹�ϐ��4��z1��(�b���h���x�^��5(-������ ���N�,�F6�#���U��t��q��熶|�hYaU�b�Y��lt�%�
���䫎��A����}.�/Z+�,�#]0��	Ǔj�4�&X73,�ÏJ��5�S���=~�O]<^ m5�rډ���wZ��>�p\k�i�H��}�D���*ByAR���$��b�Z%�H�L%%���裼�
d�wT����f���oe����(���'��;�6����ɟ��v�\�l:q�O�7H��Օc�(����T��@:ݴcm���Z��8�c�ߗ���z�����C��CFW����i~���V��7":�'�|	n�(+��*��>�l���$�[6�c㭷nB��ЄX��q�����P��xiq�{�:�D�C�5��~tu����T�
�%)�HIy��>��IԀ�Ye�}c!������`ܟ�6�����UGk��g�N:8��Y�*9}U�8��V������@ԫV�>!��T;A��tCK="�E59Ĝj��7�/z3Nc��t�e���Ę��#-ڧ����������Bd�������i%���%��wҍ�bo���|0�!�L��~�ty���t2���*��;T�I��k�{�Q^�*�O>n�+���W)�ĉޚ�W�L5�r�ӱ�7��$*��,����yw�}?
�����\D[p��%�oEa��̊���8?�>h�=�������tl�;kJ��y���v�?��Y�|�3�s��2c�D�`�ٸE��*���q&�X#�_b�%�5�@�C�� �B�!ǜVir����> +�H�0|�j
��;���@�_����A�׃]���A$���R�����_��)׈���:�2{�)B��a��۱c���A!���]d�_9���e�SU��i�j��S���\�P��Cæz<-�<��˳$ӫ�P�M�s�Â���y�F�w�O�{a5�ʮ���`+|qd2��|��HNViە�fP�Et�;�`���X��PN�Њ�SͣT&I(\v�F���h �kb�@��/
�����@�;.�a��݀45��UJ<iL��{x�����FV�p��%�/��i%�C��3^�P�`Nv׾����;7bi��1��ǵ?ߔ�~{��̎����J�t
෕܇�d4ͳ���lj�b���E���	sOR�i��li��=�yeE��GEѧ(-oX���3�¬P;H4@�髍���_�n����醳O��W?����%DC\��JׅG	��� ��3X�a�ykz�PpƬ���x ��P������ܓ��]@ɱgH��/N*�k�MQ2Ӫ������+(������>�\�����k8P=>a$��2e��E��[�����b	�L���Ņ�>�1&��?���"��i�ז����V�%���U|	:��PX@HXS3NT���~C��e��)���ڹrB���5#���<�1G�9���t8{���Ek��4k�j��Qh���RD������"��7j�6A���1 f�.W���a�_#���*���^�LZ�j�QJU�,E�.@(�O��Y���`g]*L��C��L,1�d�Ȼ�c}��p�7� >�o
A�|��T$�XL���8�\d����=��`LI�g��wE`[[d>�r�Ǭ���х�:�휜�O$:���L�	-,t��%��:tՔ(jk��>�θk4�mb�b�+3�a��K�ܬ�]	��!g^���WQ�!T���i�R6W���	%*��� !���0q<��.SIC���Ƭ�i���ɱA�8��&�^�Ds��@��\v�88H݌�K��_r��.q�����GuTLA����Rޝ���F!�̪{GP�l�e�E	�Iv���u��d�M�Oئ*{��l��1�@��䜖!�.�DX�8M+���/��z�9� �M���ځ�0���K̥�U�ߋ���2ҩ�[��&u%��-e~�<�bg<~�ۃ�R#~������ߺe~����������7�#%oƖ��YV����Я�ZrK�������H R@ ��d����������\����{�e��i��4��~���4�3�+�l����Ͻ��l61~ym��n��k��w[t�E�)���j��s�h���(}�s X!�����
��s��VjD�\%���/��Uȯ/��0���8��8��b+=)B�%iy�ߏ n�Z�ʔ[3_�bz�J>�C�y�M�;�o�Dt���j����e��⍝��Q����Z��fN���Q���XG���"���ef�������#�6���IWoߖ��0.�ny�����%^�cr��C`�**�>o_^����+x�Jɳ,�2�̬��\�3�<!�?x���K�MN�_<Ps��<��L�x��$�����9�9�^K�d@����Z���MS�b�)�Oh;��n�Rh��Z)9�,.7E�b>�2_NQ�6�n�J�)#��b�Ao�bB%�yP���s(�0g@��Tulb��15(�n�o-��}p*��.�[�H7��ߜ�S���r��Ajy�En�n��ݾ�Ɲ0���\�@S�������i���]/���P���,��V�V'RUJ2d~_��jS̍ns�����k�ts�ALc�)�-Ɠ#4y�5��فFy�\'L3���±���kU�.�aw��ě��}���N!��0z�9�^|I/_����M��{�q�Աbטp��������;S"P�L���k�GkԱZ+�g5/�<�!\���HoGV�R^�p4�OA�ϕ��B]�6D@-��rC;�^�p漋Mo�<�*�Wog�v�'���ϊ�7x��;|���
4]�]��b@�9=9���O&�����{]2�w��E�6)�!u1�P9/ֿy�/Yo����F�������$�_/߳�*�Q����K����R�6��?#Ɩ��v�1 	MG<�{��P�˰�E՞�H0��?�Z*�(�+�����yc1g�g�y�&z�O�7��X��j�C`3c��/�xVM�z֕g���1@��菼}�`!�,pO1��l��})Q�~	�|���N�!�0��ہ˜�yܕ"9T�M78���Oi�L�AS�}L��E��<P��"p��i��2�$'�]G&���πY�O߱y�|r��D�h�f��:�]�Zog�ι|As�h�p�r�y��O �骪�H���);f��&D����s!��Q�E���2��#Z"���G�a=$/�p?�3�f�FC�ej�~�'\�Q'���V��ap/�{x�r�26���
r�T�Z��D�]�{�Y�)$]����]�Eb��S�ƞyo�U�0=x�=���	��q����'K��2df&/�WD�e	i�5��ky��!�fA�H��~����	
�K���.$t��]��;�>7:]/��_�r	����"�	�J�Ve	"	9� .���}E���_�Xc첀�h8�w�M��C#�n�i@A��e��M$dڲ��N��������`���@,S!Q?�9���y~��r!���>]�T���O.S[��D�"ĝnw�7�1i�둕i�� �`�#^v�4�\�(�_�6>���t��Z�-81�\�S,v�9��4�/�Y��0_�H��~����ϻ��ݨp�rH6��a�V�a��0IEY�b�{��U�6��t�x�����<�]-��┤z+
Պ|\2DP2��[�_?��1'���;3�����q�k�0Q�gУ��kY泿��t��T}{��̄U0�3�����{�	�Fg�$���}� _fHDF�;)@��9�	"PԤ%���,�Xg�L�oYkh�=�� /%�޳C�����4|���5�.�"jM����M�#���H�C^���3��I�7l�[t�n�5��إ����ĻhمY�����`b�#���:f	���\+ˎ?� �]A�,�����~��T޳7���L�+O2B��UF�\���3������y�!��2hf������I��S{�J��d�]�t1��.$@/��}'~I�VJ8���p�
��#��LwcHb����i%@������L��ɴ�	p���� ���0 �:��DB�7~om,
�A~hz]�����3Y	Oc�Y�Ү�Ό���ը �!;
^�)G}dؑm�l�29��L�[ROrIB�� �˶�bE
���˹��r8|��tp-Fٶ=���rU�gB�������}b8�P��HI~�	PC��;�׻/�h�19b̜)\|H��A��K�A��y�!G����8��4�YP|�h$y?��X]�6<�
�������I`����+n���T���O��f��߬�n�em��N���߰Ћ��Sx.� �T���<�0p�=�}Jw�+��w7��E|c�Ã����� "�vȩ�e�J�K���[#�N�-�W5���DOk�>��5x��1��A�T�ѵ_z,W 1e�m;fQX�,�,�F<.cN@�]�w����-���f�����O�����#�M7eD��#�Y'�_(���}�\ۄ����`l{}�0<�~x��-
P��=����~��N��Yz�s�,Bl��	1:���}�k�l�N��6�?���%�|�;Wq����'������f�D�A�ӕ�������"�!�A1`��&M*�M�̗Ե����㦂���-+`��/j�;88��7��*��:G��<7\���3@]�������@\+��L�*�!h78�������CΫ�Yh�)��g�SڟbA�k)�bR�u��J�֡�w: Hyu�.Щ��k+]j���2cs6c��i�p���˥m�V�ޙս��04�/uX'�/���5(ȥ[���sb0�_5T�˅�� ���@�	��ې������	�J�ד�5_��(JMu1�}>|��	a9� {)�;=��^;@�0�f�S�*���|�k]�A��,؟�HO``�j�H6����g��o4�c��}��"�c�?zy����X�&-�7W�\����K�H���~�?��I�J��tV8�fD���Zn��"ՏL��t�_:�^
v5�g*���:5���؍��@J�aⷯ�*.Hf>�1ƑY�^ ;a� �>�7G��?!Ә�͢����&6Z�"v�Q�h^��aE`�J�}�����pQ�g��g�[��<���b�\TQ�u�RZ���$o�M����bɾSe$�r���dkX�޶���I,�[�胩ƈd���$��w���b�g��o�ss�Z�tW�;�z��%h��i[�S2M�Z�0�ηÖ����/��6 �'2��(��<�q/k����/~�|q8s/Pk4��&P�@X���Q�ǣ<�/G���-��$j��T���[� ��Q�Q�xny�O;����0��ڋ��?��h"�oy��D�&��'��� �M�����5�-zx�^�I����jk��i�(���0piחWra���oZ�-�1	��Wz?�R)��|�x3&dC^
1�]%l-0Y�*�v���3� ��e���˿��%^y.�a������%,
m�Qޜyq@�n5�Jy�+���'�%|�4�9���,�*h��z�����i�r2UPk�7�B���P�H���ꔷ��{�B"�`
��s���K[X����t+�ƠY�FWG2�ߤ����q�,����X.���2���SH�G��N{Q��{�:�z��D��SШ	�!eh`��8��1N?�
=��?Cq�=٪-���t�|�IaD6J7�ަu��}w�c�i�p@�c�ඡ��{�ܜ��
�JM�����Z@����.:_#VW�0%�st8)�UlAƷ�u5�9����s���OF�`r�F�R>�T ��k�R:��v6�H�n��Q�Zyc�d���p�m
(h�p������R���㚷k�&#���-���[�n-�@}̀I����@�C:1��	W#U֓�>k�0���� �J��XN&|ed�h�\Bu�NJ�ն�|smؓ��(�уM�+"\`X�L�Z�R���r@�7��4m��yB���z��;k�`e�8+�͒S'H��&��U^�23>����}�y��iaS�U 6�U>�V���ӥ)�ox7,�l��k��)�辻g��p�?LY����ؗ���L���ozd�rg����b>}�ہ�Y|c�L�����"F��4Ȃ����5��	vdN-XKEz�T���,��X�80!c��y6�rD������F�9�`L��Ĥu0�_�d��N�ta ��o�,&%(�Wj'�ª�>YV4|�[�0�{�r���_`��C�l���WI�����-���paR�:|��u�����e_�6$��6f���l�o�$������H��P,C)��Ms)t���,�bc�5��GV83f�C�H�t��}��'Ġ�w1�_��@��tqȗ���N8�����<��钂B0�]q�n�l]z/�7a���}S�r�R�1ML�.=,�q���?�X�Θ$*�QA��*��X���i8G�J�[hq�n��L'1)0r�2ش�Z�B.6�}$ԉ�#��]d��DY�A�Z�zp5]�=*���v׹��������"-���z����N�/��kVq�0�����7�,�܌�F��1��}�q�f��U�i�\a�5�i����ͧ��$:�n�( p�P�Z�"�ҵ�p��ح�P0�1�~=�F��T��W E�΋��v=�+�C���Q�,T�\���W�s��F��r]��"
M�u(Yk���oե��}v��:ބ�=�Y�
;6��c��ӛ� r��J>�6^7E}f�`�b��Ba|X�p�?�ҵ�O�.X�Y�ӵ�1<7��%ھ�r,�� ~����2��+�%e����B;/�9��L���[V ������.���Z�[Zu��WK��Uf2g�{d��K`?+��)�Č2B�����B���d�l}A��F0\���̴�` r�ދS�R�)��|�ǐ��o��Ls(r��˛�C �u���FW��?����S1x�#�Ͼ�ӕ�d|���܌墻Wn�� ~���֚x�h���&����J�H�]`d�E&̥�G����E��/�Bt!�/��8�;�
��gH]����IB�8M��'��kR�2@}�u<�	�|��|�-�I!qN����7r���� q�B־ۚ�:�9��/ι�����b\���x'FJ�����a�V�X;0��-���+��kv��QTR|M�EK`w(�iݫ����F ��E�)��v�<9�����	�g��]F�=�t/-���w��Xql�x�JH����\y�{N�N�~���<��Tm�m(���T�R�@M6�{F���\����$��iζ�\� (����-��ϥB��B����@��H6[�C@�Y���c�G���Y������7ځ|����~��i.��爇�)�����'�X��G���[��e}��zY"J�'&��GFA���  �j�&��D��W7�x:��廇���q���ol>�{�?�Rs����B��� ��F{��cb������b���s�'ˣD�@�[�2Xa*�t�*�0t�j�$�7�J$����xE�!��s�&�	ai�Q��Zƈ��
�m��q�B��C�;�� S��D+J��d.&��5Yd<�����s|��8A�JU8ЮŬ� �y�J#�ވX9����NN`�S~�D	�W��9��K�((oLwe@.�ua�u�gSzAD��X;iX=N6���顯���)f�����~� 7>G2L�;z�ӧ.'����sZ�(P��jp�����ݽ��k�hS��#�Q}5�j>w�q��܅g.��W�����[q��h�NG�3�ўOv�Q� �p*%�}&\6R�e�n���*�����7��`C顎q��ڶ-��K�=B0S�\�m���'��v�6tȧP�:�Z�]��qu�F�"E�|d�$�����DK��05�K)yr����	�����(�?ȷ�S
���m2�Y=h���&c�D���m� ҍ�v��ӑ_]��uz�\�����\�uW��C� �d��8�A����H"i��_��#�m�g� lIU/-w��r����H��=���"f�b���A����ϻ�4l sr�x57��� H>(�V=�P�5�L!䤗�� ZY���U޿��ڼTvLoX���% ��M���Wg�������+�_� ���-,�U�y!>f��G�N.@wu�A����8���,ch٘�{�9�D��\���_������p�7u��1�[[{)���Ĭ��Kf 6�L�=�p\��|�,'gt�[�^�Ri�E�k�-����5��$E^Aq>�H��&�`����7�� �nȐ�9`H�T]i+T�{�� 	`k�ҍG�K!���-�2�ײ$�Eڞu�T�� �;Ab�JiQ���*��E;��L]���O�1A�kS�U���= 
&Յ]���n�(����U�]���u�R��F�ۜv�8 XmN�m�����<f�)0�����sL�S�����K�������\h���V^1�T����F}���?�����F�F���B:d�8�����na4�� 
V�+~%eT����k]m�Lo�Gi����nP���� ��u����*�������3XfK�*ޗ�c}#������7��G�7��r�������0.��P�9�6��W��;a���+�Fĺ\w�#���7�#d>��7�!�(�h�h�<�oc���ݦ�შ�ukk��1h� 欳�"�|�Sn�Z9��q�h�q����-eY���5������$�T��h3s���n=��P�Ɣ-�R�wG��m�E������I03�z�(��f[C���E�`=�e�n�ɴ�3e� �O���~�Fp�PB����^�r��7F�.�O�|ū�5,nZ��,���UaEI	o�K��?ma��H�T�����K���:,��K�dnx)&�sc��]E�i �s)|q2^DF�G���P��a�#���L\�g[�>�E��l_�\$��Ƈ�'���BA��U�h޴F��A��*{��w3�>E[�O�&�{�a�JQ��0D��٦b�YQD+w�v��9b)�&T(�\v��� ��ś#u�b��μ�Ԓ |t���X�7�*^��� �#����A6�b$W��o��[��Ű.�@]ukC��ө����y���@V��_�=�|GUK���f��?f%���~�L�v;*@���M�1RQu1�1�d�u
fº���w?��X�҃\�Ւ^�&��s��*�٣��۽8aH�2�	*�����ހ�.�m��P(�|w�$go�8y�ؔC��2tD�ܮ�(O��O��� ��%͖���$O9���hD�<{�a�v�N���9��{Xh�yz��i�c~�\Ci��-�J�w�F]�K0�8�·�#D�r/�>��"���t�܄�D����}"�%)s�h�#�����V߃����P�躸m�4����]®�/F�O��4��@��u("��$l9��?(��!����y�Q�Egi��Dz�졾D?#�enb:�FߥZ>yPi�d��,pEu��Jw� �x�IzX6����vܧ����n��F������a7�o��7��|b�Bcx�A{9+���?Qh�Z���{��>9�����.2�
;+��BKJ2`����S��\�1_'8��8��e׶��A�=�`V���Y�#D�(k@�fB�V*q�{�@y���b�ź)��<�(&�*�AV�����}��`���H���Y��oʅ$膇��7{/������(&$+�ދ���b.w�а��u�r�%J~ٮ�5NgDЩ����pHr��B��N����<�:]-�Ļ3�7�G<������8�ū�-* {��J"�D�Og�ˣ���A���T���o:�����K�P$�����$�:�ႃ�����/���z@���y�f�ݦjyS��\���d&˸N,��K�圯�������U�<K��y��CY�Q��L0 '���`���1r̀�0�[��>Qz��rg���B�6����c~�qU�c7q��(���괿-	Y��������rX�����I�sN�p짿�3�{u�]Y�J#�q�1/~V��H��І"��@����`�����0�W[�L�_*��e�-�-���*�5��ŦL�U[$Ҧ�*��h{����"���3Zo
�,J��v��hǥ&�i�"p����CL���q�E��@��U,u���; ��.�lkQ�`d��4,Q�@����Ӳ]����Iy
�E�ƱiU_�N��H�ćc�	7�L��2�7�V!�`�� Uǡz�Lܿ�B�g����?��Fz٫K���^0��i?%�P�,i��ԣ�D���)/�����*��2��#��@t< ��b���?�@�A�X�L�O	Ǎ��Bz��B7���.fr�Dx��LH��>mt�1N�/�2(t�vw�Z�NA�(�ݝD(*����<���� YaU����i�g�~�w�>$A3���*֪�V��۶�eFKXn�{a�/*�l��:���jo�?i򽗘������锔c�WMԪ�d��z�/$THg��<���"�^$�p�C>.�'$�c�Q��!�fv���ɪM���L�H.����-��*U�(�����R/�ƺ��g���|���*n^p��R'"�L�M@$)E��L��U���QJ� � xe1���,Q����!�XA�]����u���Ѻ��v��A9�+mY�KAZ��`���b_C�'<�rT\�!�񺪃Z���j�w;�S�Iv���Q�!&�����V��1YU��o�]U��M݋���k�KH<�n����T(����	2
���<��Z�_�j��Փ)����1�ZH����:c�=$t�K�L�������;*��I)��^���ɟ�Yƍ�6e�`��W���^�)�R���/<z�qE�j"��6����5�V��X�^߯�Ǡv05����g�f[-n<��#�Uq����c�z�p������y@1RR��q��q��u��Y��� r��G���Ll��]��c��N�}�Fmc�9*>��%���(J����:��+�5���b4� �����E��`j~�kvt�'F;)?��?�뎷o���q�0��h�nCr�I>�)7��ʴqR�W�X^���0Z�����0Y`5��ψG�� !�� ��*-ϋ�l�;�>����X����~;Å3�~W�W�d�#�֮p��r�@�{\�_�����=��Lw\�~�D"z^��`RH�\;iwХK
�Q|�7�L�zLX|o��T�s���F�'��4q�x�k#�YRt��?}�d��B�e>�bu,��ټ�{<�a(]9;�[���1:�q��\�Im�y���pT��&]H}�-�
�]q�,���q!^x�Z����1;N�3Y��=�F[���jg��Y�:ã���  Z�W��(�R�أW��<!�/>~`��~(Գ8�T
�>�1�mx��Gfu6u����1�n��	*SBN/VK����G+���S��D]2ǯ�2^)�L�6��(�gDJ�a�y��9QH9Nn��C�oGz��w�={�ט�vմ �jU25��t��9�_��<�C��@����7܎Ee��-�3���u�UvuD?�Q��@X��ɡ' �D��^�?�Az�����$$_�a�:�<%O5Y��{���ә���˟�-� 2Ji�E[���m#�@����~RI��{r�$CH.����hdP0T�X�R��#=B��2�a�mz�!hFG�<\)��ҷ�|jy���K�`V�o���Ĕ#�'ĢK�������5 ����ٟ�o��Ny���D�Ȑ٩�W�GG��x{bO�d[/�z�#GN���_�W������ci��|_ɪ�\���y�R�ӯ�kʼ��$���u�ZE�PJ�Y�3.����k��W�|"�g�$����ԍt+m��p!M�t�։�t��t�#��R� _	��,�i�4q'/I����� ��o�I�3�3�
|��|���=ӼȚ�te����"�0���US��r;�f,Lag�8������\VM����W�M�/8�c�T6�4��xO��Ȩ�;*������1'���<[g�h��(.9���o>sʦ0[.b[!{�%��^�.�vyg٣��>�>���z�ݽ��>�2H��I�9i�?~�7gAI��
�[��}�\{��$]3#~�m�/z��H����M�P8�ʭ2I0�)R����������ϹPл�����e�8΢�y�h�S��
Kq?�*4X/O:�m=5E��P��(��+������;i��R���ȓd�]B���hY,�&C�׊���X#ZUI#��\��O�&5.�D��Ux���0�Ӛ�4��d�w}0�pX�$�!rf�~���+�����[&϶Qo��\����*�l���E9aɹ�b\��o&ό�����Py|Ө�i����"?	���q�l�X$Ч(�(�(l�̸���Ѩ�7��5�۠i�Ze��Y �l�Y�~.���������Qf(VN݄��,���U��j�������>?�^)�L��%��=A�l��b��y�&i�&���]I�f��,��y�������$ח2P���}1F�ꖲ�Z�,�k��ñ���S��Y���m]ؾ��!��]��è�Q���њ�������'V�<���_��H�?큭|��]I���g"6�6-{������z�_
�JM�KT�}ǐ�P������}/�	�,��M��K�p�A>�!��]�_��܉d�����ao�ء���ɪ����|�K֛5FEAicbJ���*�ll �3%��Ͷ�yՇ����W��!7ì9n[�Pզ}x�w�J�jg�A��)D)��:qP��q�L�-Y�'�%��ꁮ��߲�n��b�IL�	]T�]��ܖ|�8>"I�r֓U�b+��
C3�l�Fe�ʎ��'���Ϩ���D��*p���L��P�b� ELdz8�$�7!�x���7�1�})���>?�C6�B���E�ﲚ�T~'c����hcؿV GML(�:0���/q������j�ۛq�9���O�$[8��X�7rfܚ����61�]���S�:� �Ⱄ�#HG��cU���Z�5�V�O~?&��}g8�v�
d������+���8g�|�%X����cF[_�z\�%�YԎc6��v�.���8Rh`�7~�s<��7���Z��iPM*z�~r�մ�Do�d��sXi�ݨ�{&�M��n
Ў�W ��n	o��|��Ю�A	�b=���N������"�Y�_��Q��)��Yܖ�aYy��Vc}* |�A�ky{��i��������bP�k�*���
�w�~ ?X%_	���G�R\+Ǣ�@:,_�I[vP%c��#�Ƽ�2��߾�9q��G�������9�! ,#a˸J�Q���X>i��P'WʐT�0�W��%��G��n��8�o� �V�]j!M�]DV�q�R�)s^aQ+���M�*�H�j��U$M�媢9�@!Oq�i�T��gFbapK����Eͣ��4���b2Wy;g����@�5�d��d%%	�(/��Ȳ���4�<)ԣ�2m4B���C�1����� �v����w���>B���X��t
b��a���i �f��� ��o��e1��7���
�e230� �{�`�I��V<�k0����ݮo[��n��}=��q�ާl��v���g���U� ���c��c�	w(�Y��oa���%�����ġ����8�������-.
����m�	
t���N�*�+�]����9Q��v��x�'%T½��b�X�{�J	�ۜ.v}��(��@�%�i�&-{���tl�~:�ZH���pO�(��w�!S
R�47.�Η�C�cs�@���{�����
�y������!LP:Tx%�	�fsy�?"��t �q��t�?B��9����1��D�8W|Q�j��T���mi�41�����Ǖ��,r5�aD�P�ɛD^�߹>�<����V��ɴ4��D:���D9\F�"F	O�H9}}���:̠�"#u�$Y����؆PK���.���ӊ�U9�8�L��/ֈ8�y�V$���z���~�Ʒ��4=�M��� ��$b5�{&y����e;z� �ż>Fv3,@��7���>���zJq.�
4�k��\�.T`�� ��k��;����z�ٙ%�Q�`�ش�h:Z����ご4?�%�qԗ�1���Π^usv����=��}2`7�?�DTB6G�ٝ��R�S���T.�����4�0g����q��H2����P]��2�^��]�)�%%^k㵵�e�<���-��MF-�3����g泝1W���z��B(�V�v.]lx�X'����;��	A /T�g=ǻ"�s�PbD
G�-?�?�u�w�Hq��z���R��#����Л�r�Xpi�����
� yO?�&2��~W�;{x���'��)�L��k��=ũ�~c)p/	-bM��B���K��أ//-��]�������²%���tkۥ4��d�)�̆�. @���]��}z���:,�c�,	�ѣ�mj��ch��+���3;�M���N<����@n�Mƪ��?'Z���N��C��{���W���/�qb����}�&��Q�g��[��
�q
�GW�,�.��=��h�=�#�8���|u�a�Vsw�0%>���haKGgۡi�H7|rx�+p�2C�U�к�2�3��J�)�%#+���Q&]���l燳��UR"o(ﴐ�.�Nׇ�N{ ���T��nep���g|��� ��7A�'��7�C�9y��䗿�L��������83Ɔ�ET=�I�}r�Qј�i�hl�G��x,��c�����7�(�4Y����SO��nh����M�e,a$F�!"1x5�c�"��w�����,M����j���c�誒f�	5]�����������P�,�򁒖�z!|��,1��w!�	)[�d#`pq)��C�^��w/h��dy�3?u�Cp�K�)n�1Y~woB������^%��tG�����b�@���fM�r~>
*P���UА�S���eҜ �����F2�0��H0��!�Ѧ�7�o�4	E���~� �б���_N���$$�����ۭ���M�6�w�K��3(����)�>4�.̋�,�`���)NQg��BB�ۢ�)��ٮ�_���u���
��?��"�#��=�U@���bdυg��g������������WE®_��Kҭ͌e`�0m��i@0�j�rJ)�t��v(���F�H������j�� `��n��~����2Bv*�$���㕯��u�'p N�IS �gK�ܖ7�1��<��m����lQ��F��̣\���BqP�>�K�ׯ���=e�5i�ںn��g;�FeYpy��WV���v%h�:��#�0�ե�,�;rb�UhP�R��^��
���uN��3�Y���8��J�a׌Jº�x)a:(�^�)�^ƿ.�GF�	�!5�k��ڗ��y�t����F(�*b+��sS����h')��䳄~���pA��q���c����g���[�f)B��C��l5�S�1���-��c���JP�� ��KZ%$s,>!Ɔ7�1U&�fp~�ޞ%ǩV9(�wGzF�޻t������QGC���9{�E�e��Rp��t�~�g�so⟱��GC��������)'�s�`?�ͬ�s#)\��T���]��!N�`�NO`5��݋��RY�p���Hh	X������b��a��/��q�G��jpj^�(�$�#)E�l1��`� ��݉�<�Y�/�������Q޺���f�+�ue��ቒ¾��N���⌵L��*�B�%'Z���Y��n�^�?�}󟇙��Fzc�g�_�[J2� o��.�E�
8شE�xY�x�GՐ���hg����,[�y~���+�Mt��4�`]VP�\9��F��;g�4��OOW�X>�{mV<�~�Z�X���8L�1�	D�D������|"{]��׻�3�f�H�M��<5���e)�W��噈�i���'�V��$4fu�cВ���,AP[���΀���Q�Z�!�� X���=�[*�Mb5|y��z$F����EZ,,�E�i9d�Z���Q'#ź�K��=��~�b�{Ȕ��]P�Y�Tg9��4D��_2�%&��AM�T��1C�zI��5��Z�����:
wM�{�9�;���o��v�Ӱ=\zGe�4F7�M�/��&)w�*w������H>�.�V~Tj�+cw�<�i$�r�����_�P�s���� ʄ'8�a�bs�]%�fZ�1����y�q���1�'CbO�N;O�~^1�X|`�m0)�e&������6�׿/���B�~�VY���_w 5�4���8���}��O\�����A|�Pf����9���X��>H41ʀ��B����ݮ�;�L��?V��7�=�{��F�ŋ���nM��t�a���W��v��r����.-�zx�[Qh.{���:h����7��r�99yb�<kQ�����(�L?��#�p/�ö�U����؈[(�̸RYG�θ���h~W��tm޿�Y̽���!1� 8�-"�p��gʶS#��U�UV�a�a�M������c��Z����@�"��c̹<��=s3������N#q�wR�-uE,�57�%z���J��Ez^���4d�]�\��E!w�I�y�3?1�M�Э/��V�6�[a���U��gg�݋}o.2�V�6��Q+(��~
��D��z؅�W�}�k�
�����y�Hp'��x(���n��aN-�%�>�	ubI��������� t�8v�44�p��	��l���ZO��W!����b
�u0循�[YE�#lH�T�ݢ�o.�;M�%������N�6�7u��r����r/r��
)��0Xh�̣��y�A�]�����
C��ö�%�QO|�Z���}�!m��+C��7�nv�/E��ZN��{��ҷ;�dY���6�<4t�!�o����i�_3N�G3	x"_���aXJ4�)�K?����@�KM �9�uB��҉g��zSnC�_���y�r��	���Q��BZ�y�hN���x��Exn>�:�8���A�[l��wUw�ɵ��ǧ� ��v1jDyhP�ޚB�x.R/F���~�[
CV^��#mt�s+X�;2��]%�<TdJ���>+������ғ��u�;����2�ۿ�FPxXi��d��s*w�s�s$���M���Ζx��Z=��W���ǰA!n���P�[�$���v{xR]�iu��{�>��i��l�蠗��v6TE��b	���?�N�����}g�y��'�4!	7d�ʝ�-�齒�o(i/(�ft!BP�@�})��5���q*{�����$MAp�8h٩[�{�O	h���T�f4����3;j�t�����gv��4����C@���n�t�<��X��3ag�9���Y�X�dYPlH�"l*eH5剣�Ÿ򱓫TY[�'���%���N�+����P���n��+`���B���[prG������6��b�0b��B�p���$O4�N��=0�S������Sc�������]�_���I�mZo�+�\c(�R�'W����>;EB�U���Z�O���`\��(�y%���Y)���(kؽ!3����E`�/Wd�9�E�gڇ,����3��7�Kc��=��jB'���MC?	Ǥ�$)���|��b4��p ͝�w�t]p��� �Z7��_@�e{¯Ǆ�aU �<L�����㶨N�r�'#qJg�x�3ݲ���ʟ�m� �1l|l�:��' �4�a�}Ā�RsHCm}XK�av	��[�E�[Knp7ӿ�GU':֚�t�k]d�7�� ����*�p ;8*��ɖ�E"$�G	f��'� o�<�H4�F+���#r���?HM�\��b�A�m+��@g�I���D�e.��.�#��Z^���p\��Yº��Z��Ɖ�,"�>�["3Cf�*[֎�X�ˢ҉�F�e���
�;�K9����t�4Q�(�����u�u'me �/y���׽���cv�Ko�����SIv��hc���R��Z�>yGjnB�����&���S!�}Ԝ��@��YU�8�뾇j-��7h�~��Re�誇b�g]���\nW���	���?�+��A7�k����%#�ԇ|�T�>�=)9�}�7�I"/R9.�kE�0B��	i<��P�s�p-�`%�2�a�p�a�J�y���D��3���.9�H6���&yK��
c��z�a���:��Z =OD0��n��2�h��m���O�Zi�t�[��ϋGֿ��%~P��L�)ϊ��l��!�95�;���߸��[�Č^7��C������vp���4��P���Z���)�C�2UJS�c�9
��K�����f����JJ|�?����a�ҏ��ݗ��x9bwL!�˿����({���o��G��	K8ȗ��%��Z���F��,��r*�U���,*=�gךּ#���Ku��1��.��=؇��8ǩ�ԕ�>ؾ��vD�3��s#4��]{�U�I
}�
��I�b��>7���3 ��B�n$AA� ���(�̳���U"�d�;v�8��T�ws��ӵ�/�yՄ�"��G�H�Q\���#�]�6b|�eXk������P�%s%�X��m��~d���CWҳ�Ɍ��eY?�?
D��D�h|�5�WcC��+,�!ܖxS�J#�p��t��T�;���s�e��Gu����d��>F���Q���w4��?���WΖ��b���?�:���|J����{ ���_��:8��X�#�v���b>��y �O[��\�S^���x}&��v����FY�Do�M�V�ÊX�x�jܠz8��6��!$��&�I�\2f/����vKK�4*5Dm� ������H*��u�m����^g̜Y�8��#��!��"�=l�J%/�{�ឲ��=M�6)��w^�n�S�JF"�y"![�K<���x��Xh�vu4���5��Z$�Z�E:�l��IwL�N0�W����%u��>�%~.=�0P�3�ʸ�AV0[nD�AʹP�p�`��6�l��RL�̲���B�\�G��OTl%Z��&5�^���t@X�Z;�G�>{0����M����r�Y �a�Q(�TK��З, \����,*N�_��?�U���j�sǰ��NK�S���E���(Vl���p��D$���^�� ���j����WW"��
,� �~�Y'���z7NAr��
��!S�C�I�:�1;�jԯ����n���P�
`i��	E�tL���V{h�`�6ceZ���e^�]����vG샜8����}~� ���&�-B�
J��P0��Kы�h��
G��<_4Yϵw\��8p�뎖HH���@��OY�� 
ūK�����#X��:%���������p��m4y��o�F�Q`�qtt���Wu���k���@S,����)>��/ y�xs�í�w�6�i�t�U��_��r p��^)�;#�\J��
@������>�B��\`��w;��P,s�Mz�W���*";,u'��:�q�O�-����ʞ�7#��q.�4:�6�;c���PX'��`�-���Y{�P@�~A�IO�~c问ݵ
�,�� >���9)*�e묡5��*=~�q�H_�M�5�
gVzmVs�I��tH�7�9r�e�����͟gr姸�ye��G-�݀Ļ�u6˲��C�E��)9Q��GR�rө���]�@C����5����P1ĦmCP�↦�c�����n9���45kӉ~��������y�Kf�6�t����t����4��֥2�<&��(ز���>���?;��-���oH>(���3�u���#�N,'�����t9�4L�.�1��2��M@���~�G�>�Q�S��4�s��.XɄ��ڞ�U@�s�^��L0�u'�j3Y�!���I�W�dir��lפFK2(���������Rv,5��G��7�����R��!�"4�zf���0���\&WʽN��S������x�0r)��>*�2��mb�����Q �6��p�U����I�#ã��DL�����{�0�x�3�W8��;�W���m��.�_64-cx�X�w�M숉i�H�4�PsAb�;D�3����]���5Q(ٰ[�jh�n,�f~� ����K���nt�a�e�`@���h� G��-�5�a~Rf����N�DX(9W��<D�u��W%!��t��)�D�5f	ԝ��dfv&�$���U2��?)�����(�yn����{�
}��KBi5�Q��hU�M�������ϿH��e���a0�a�o2�[�{V�g�?d.��/[_��^��tD""�&�ofzݔ"fD2�YF�΍���iO-:O��B�MDl���B����o���͐WĂ�ɤ�"K��1�@"�z6���VE@$���{�g�?����s��7n�ƫ[�в��*C�g��V���m g�����#��vʥI|��-��;�&�q�5���^���UbZ�?^ �\�Ls� ,0����⼓����_�x
9��ݿ KP�����Y/�X��x8_�egF���E�ٖ�9p��9�Ǎ��i��_�g�kS��y=�~�Օ�y��	s�m�42�ϼ����E�%�Xs"��\J '|��\]�`�i[&�Z��'���۴*#D�H���;�׫���Zn�i�$o�t�Ǎ�G����\&^}�y��`�J�QlK4�,�R	�G�M�VK+��F��O]�2X�\�$q�Ea��
��ܧp�?�3K&�V}9�>T�c�(~yຍ���V w����������L������],T�p��r:n�vv��o5n4��m �-�(��̙��/���;�o��g����3o��X�G�j��\��`��}R�#tE�|\�p�� ���+"�yWTw�Wn�­)%+;�UN�vܲ
H�!Re+eP�u[��]�����:�SW�Ĭ��~���&�M������#�{^�Q����%m��h�&���$f���(��4�-��0k�h. �M�s�y�;�f�y�ptq��!JMjM/VT;����#Ja���N���i�$4�#��b��k�*+х�EO�Q��Q$)�<B��&5�T՝&�R�rAW6�'�.FS��7�G����^밑� )��tJ�B�gP���n�h� ��a(�=�Ӯ�YWA�u2lq�Ҝ�y��pd� Q�!;�e��2�t�P3�	�O��5y�DI�p���N9w�(VvE��?�����?]]-�A��n�?�������hu���:����ܑ��.{� ��DLo�	p9�I&ɘ������e�P�87I>�}W�<R���;K&E������P�h��͒1Nt[Gb���5�f%����"��\bB�7��?]]ϱm4ɟ:Y&'0X���ȶ1��X�Փk�t+��*�j������~�4I�>S㻙�����+�k\K��Lk+�N��]1XGW^�݄_�0���0u��FXA��;�{va0/�=�/3T�����(*���lC�b�"qqz��VS�<���ߴS%���iܗ
4FJ9��*:�R�T\�>�|��]v�툁c&!�!��HE�X���[�*���d|w�Pf�-�[Ǹ��;'�ƨ����.A¸�����j��˿�0�?﷾�v{���|�X� t;� ҜW��B0`��J+'���w4o�	�Ї4���zusm��	~Eʄ� ���t��|$��:�xE�����v�4��ڌT۾����Di�����z?��bI6|�&L*���'3g ��� �*�Z�LY!�w��I52!��	b��7S��\�b�I�8�d�`U�0Sզa�o�ʲ�q���#S�<K�FȷV��^<���E{������E���D�+��X5^����X������!B��S�A�sx�_����+n�;�1��q������@�m��bv6�7A���T6��t�&#�^`�A�Um�M�*�R����7q��e��U�#��?O,�{g-��������oin�����Q��R��0%��֢���׭����
~��y��	��m�;f��Æ�����B�{�ZXy�5�JUX��R�6#8��Н�%=Mr@��[�����4�i���Ff4~t�̂ٱ�,��4��eN�:]C���b�ŊQ2��
������ ^��Xyr�m��g��{d8�Cp��k<3�X"AL���rv�G��/���|؂���(��H���΃0syF�}��ˎR�&�|��ߧ1/�{+U�T0��v��yA�i�i���S��o�����c�JmLy� @<�a�s�BgT��ec��R���M�C]�x�,Lo���rm�����@�l� �7��U�k`�L�B�ާ>"��JSs_���mƾ%mW�������7B�
�Z ��7:�ټYqM���[J��_���h6�����.r�'��Z&kߝ�~Ĭv�'���!����m��[�vF�s/*�p�t+ID���8rӞ���ʔ��H�H�����[���3�1��1ʵ2��nz<G<��B?ܙ˹)o����8�x�\��*c����Se�����x���S�y&�����/����п��i?�`t¹%#��J�m?�����j3����r�@�C�eѽ���s��S�a|�<�5�ʓQ�O
t���$�p�<���:�+�iβ���o1�w�p~S���}��^[r�d6ĉr�=���<ʈ9�r�mDT���RQp��4+;�����_e.��<U��vƍ
����	h����}y.��v3E����	�>j�D |¼D�ӂ)w[�m,��d爐]W&3��G�N��܁���ZY�*;����Q�:J�a+}r���F�d:��������,���.��@��i=Y`/zW��� �BU�h��{��.{*�%(�t����<���ۺ���!ڐtrU��K��A5�}��nH�&L��:Ȧ���Z���}k��o�~9 +N|:�x`_د����a���9�ohk.7�AHa7���N�>����y�rc�_���\.����X1NRb�$��vZg:L����Zb�W�Ty���G�`��7�Fp	N��uQL��y�����Y#��g�,F=��^� gՠY�Z�`�>�r��̔�+�����A07KP=�������h�-BF�\�Cyu������d�Խ75F;�� ݗ�"��o�{��h%����#�lMX]�L <���6�P�أ/�̓��\�C���-����2��R��r�-��z�f�V��A��4o����b�He<6F���vI�}�ΕJ}�qA�h鐺X��U�9�r�?
@o��:�T1.�[�H7G��cZ"m�KE���x[�Pfe���1e�������];��� Pc}q�]]~h��V�GN<�e� �������$�E�K�����W4��R	i����(��:/%`L��-$�����6O�3C��Y��! a.'�h����6��:��[ \�΅���l�v1��LJ�[�'Q��Q��6�X4k���1�����L*�6�L��Q��ha��lumr���%�cA����+֛�k��tٱM`*����*����ȩls4���E'�4�(���ꅎG��]�-N=�����*̩=w�{4��gG/h*�y;1���>7p�<X���|A#N�TS4e��u:n�q��Mo�v�Pɸo���e~�:K�F��Ǩ2Ӆ�CS�_���h#-�,3�6������Q��AӰ��b�ҹ�d� ��v ś���"�}U�{���3��7���ы�����{� f�_s_A�o�}�At�qqR�k�Wy�	D=Pҙ=l}^-��~�d�ͽ�f�O"�J�6Jy^%�I���v�C�W��aC��FƋ�߃�C{�l) �n����X5
�U��݋�:�V�~*�|R1%�$n���	�3z�3��X[�i�|q"�ޏ�	O"T��s��n���F����%�"c�L�J�6A~!K��ӌ���.B��`�C���@0mU�����BT'�Բ�I�/k�Ǹe��@c��3��]������(=�,����r�e����Yed�0	���Y�C�΃rF�`�a=翢S��2�B4)B��]:s$Eag�鍌@���Z1�����TYW\���`�`���+>�i�v�2�S���� �C��M��>^� �qļ��[)_}��K$����&=�-�
NӔ�c~�<	KԊ�'��e��;q4�k˪�N�� ���ښC��mn	�Kvpc�V�
�*���2����K�,�G�P#J>e�h>KWU_�?��f���ۜq��n��U34� �إ�
o�A2/�=�+}_t[��c��s9Y��)�wy�v
f3͑[K�M^��d1�F�7������-+X<��D�X�EGVZ��!2���6��Bf�#��Hҝ�l��N��i� &��c��m�\a��c+Q�P��3(2&$�m�D�4p�0.�j��D��{��Q1�ѩ<�܌)�MS��Ԑ/�:8.+��*^3p���B���?:V��k¿u�t�(s���C��ڶ$�׾6��@���ϣh|��g'�dȾ����Cja�d���)�R��{�cA��SAR�4i�XS-E�v&�N.;"b2��v�����ݢ�e稆�p:��[W�=x����$6�؂e@�&�.I�҃R����1�G�7�O�Ą��̌7���h�w�5�௝�\�Y��s��-'sK5"�@�Q�!@�Ң�̦��7�,�+_@Z8�":�7�P.��>���H\�?8ڏ5�eO2�0BQ�����L~<c��M<�v9�C@ľִ2s��`�<����M���Q�!��I���W��������x��L^��& �|u����U푆A!�ڑ�׹x�,:��:x5V�����fy��s/��²���_F�S
O������+�~���ѫ��k�S��/���(�o���葊
4@tJ��S����7Yg�b{u1�]׋S"bc��U��h�M&+���dL��G� S<���;e��6Pth�FN�R�rpm������LW�a�O*"#������s���8�h9LEZGb�إA�i�K�7,��B�R�J�V�O����z��5C7��H���P3���be��@��(j`+����B�CTE��*�Ly��]���6���b��X�p2x]�%�V�]_��t�Kͣo_��>�BƾO��$�������i�'����!�3~�|�@�2�!h�	��Q���N��^�;��vؘ�6�z��C��AH�{������<Z�+y���u�^<�~���<`�!��,���1�H�hV�8X��Di`��=q��9>Z&1�t�I2:��E��-�Ƣ�/�"�a3K�O=[Hz��P?���j�>��<�c�i{oK��?9�&"kE8L�0,7)���bS3�ȳh�T�"r�7:�ۂ�C�0�&��:�j�b
?Hl�t����Lr�I5Acd��T�I�mY����Z-p� ��K�2��NG�=N�D���p�34�}��ܪ�Nƿ܍Mn�]~q����sh��-���R�n|�N�"�_�f�����GK ����:�K�>�����O���h�C�N������,Թ.3G���?<�b
Hx܃�y!Q3��)&8�H�8g��I�#��c��B�ͅ���N:oA����;��Cn ��pJh���?WF#���"Y����=�9Em�ܜH�Ψ��)XeEL����2�2�G��a���L�F������/4R#�kD�5�q�n� �O>̷|��_���޷�ˎ^0V8(�sl/r,-��م�f/�ќ��A5���ڠM�j:QK���-qd��?nҗT-�T+������(h��ǡҦ��x�����6�zyv�>G�&Z�)���>㌌N�t��s�@�k|��	��u+Ѷ����(��<��~�Y[y�C>h�v"�&��SV\��9kπ�u�R#�7����A�hݸQk�T�|�(�*|D#�/���{����Ġy�����?�z�(�HRqs���_�ݺ����Ѻٸ������o�sO��/Qi:���8���_�6��,��w*�c"���]o�}���g����\�\f�s�k��p>Xo!�$=�Y�K��Oԟ�3�r�;�NF4Te��������[�3��r ���x����wS�&=�ϯ���Ԕ�G�Jin�����:��������>ME>��1e
k�I�KK����`e��%��i�)���$�.���a��!K��Q���t���V��Nb�T���rkM�GGd�`��1xR<�W&̮O�����V�!���O䓘���i�������k�e���85����0TU��p;������'CYӪWV��ol��c�'�����8��������k9~̓s��]�h�r��ݻ)P��@�����9��kC��xc-� ���hsC���s�4h �9�B��q�����8]���$��y�x��>$�v8W�Md������1o3D&$n��!�=7�����&���k\]�Oj�r� ��su����exYq{W�T.#-��<�����6��TEv�wF�U��W�w7��^�n�����삜 ��uW;�;����`��M	�5	��Q��M�ͻF�a-�˸�"G��G �P]l̺�z��9�=��^�;�q�;��b�����e�1z�%�6�I�����r�q?O��M��8����)3���בaJ�=�Gp�`�Kh{���l`�>>2D����?�{[?Vq����mg�ud"	��E!�r�'�R#uk�Ƕ㬵j����t�&��I�I�8/�,�h��{�xm͑R�%��x�K1X�g��a�=~�!��?� #�"�T�9���m��Ql�����x�%~W^ޙ^@3g>UC*�q�W�ɻ�V��-�e�m!�~���s�t0괝��F q����� 	�ۅH�P�Y�y��{��j�oy{��)��I�OaY�뿢	Jz,ı�hE�W�YV�1
3$KQH�!F�ʏ���%����ܵ���ۇ�C�h��3q��ӧ^�p���<(�|
���Cۈ��#�I�&U�k���>:*��gT�S����ܐ:M���.�hڸ�u4�^��(�p��H�4jΚ���!9Ao�Q�'�PZ{Pb��1���b���c_Ր��H��'x��TI^
N�� �+��n�L�y��4����;�l'�5�%��gzpF�m��qGp{.�
��71(H�[��Қ}E[��ʂ^����<X�s8=�o��̗��{z9��n�!�O�o�a�絷�´�73�� r=�q��ݠ((��}�_�d'sc&�� zN����*E����#��k	Ŭ5Y�_�w�^[�����鍡;ExP oB2�a�rm��&����(�BbԽ��'��!�\#Er��j7鮁���y�v���bնzK��igw�f�@�{8����:]��΃p��S#��G=��	43Z��=د���zf�VS�D
�X~r�c-���d�Cjlۅ���Ss��
������� 0��|���m��j.ˑ>H��;�f�"!D�o%7�e�E:�|�y���J6�j���X6c�f�wU���n��t��3Kg	��i\�h�p[������)�>%8)!���o�X�Ti%���T�ʕ�6��2���!\+�Γ��pڥ(�F��-�1Q���,�a�i��8���g��Nְ&�U3�iy���+aR��.A����|���vv�e\�nO���Zߛ��������9�6q%s����(*�L�ܭT\Y/�wA (Pk�_B&yv���ù;h=��[[�Boۍ��2D���d�~;w�����n��g.*���fX�'���Ϩ#��i��+���h�����^4�p�-nkz�|�,��1&�Ҵ�VF���MeK��4���R�-"��P��a�t�׳��R�<G1^����.�9X�H{T��cփ���NM}�4�T�<;�$�wr����sN�Lk\���B�Ppf��>@P��M[KC)�'�ql��!��ײs�w;3�j�k�U��l����PD��Z�v��<� �Q��$/�>�&�����a�������}:y��]�J��c�?���Ljd��[�#��+j������cZ���� ��r�dy'��t�g��D[~yJg���N�^h�yCߛ�_9�B�����Ԣ��_��.?G�f7$w�����n�a�~<(X����B������}͉���a�3k��C�I�~=���I#j��Ho~?�b��?p���%�o\�e��A��<`Ɵ��̐���yx�����2�
�O4���o�a0ػ�@��/y�=,�
@+r}烇?825Pp���$�c�a�v?:��V���Vr>!�;$���[�����cɰ�h߸dq��*x�A{���С{��=Mg������k -{o����me	H�[O�2G�m�b]�m�}W�'��c�,�@	����糺R��тt���k��3�F_Of�Y*mvO㬒�z��G���������W�¼��U�m'n��>7%Yt&Ӄ2����'�o�K�j�Z��u~�]&�������r~|�&�Wڴ���cB2�s�����T&�ޞ�Hʚ�aYq��Qm������5��5�����R�{-SS���Z��a����w�
�����Z����u��M�W�<�Ģp�ا�ҫ��	�&���]���d�WEfo=�'5S3�u=�N�|?wpQ��飏�Y�GC�|�em�P�F�5"�V�4J���m�R�V�<�ӦX�C|��ć� <�rj�	�Y����<����3���o#����뛦P)]8����^�2��	V����yl0��5*t]���'���r��\Y��<�6ߜK��%��beA'�1�a�J!O��R�+C��Ext��ˏ"i#��.�@��m�����P���8Vi
�U^c��V�+���C�nm��ָ:�_q�"2�3�"ڗ���jr(����^PUw'�-�\Z^�p�%0:{�����}|���P��(|�.4a<�6�UFH��ٌi<tH�F�JW�;��_�F+�u�^�r?�a�C��ن�����?��(�ћsK,����>�s���g���@�kӏ�Y�3�{�_!a3�ҘW�8�==x�>��Rt���q���:�[�ғtґ��"�Axc��Y�~�Wꅸ���dد{�,�'�jPcm�9C|���냋�ߚ�LpT�hu#_����]�/b���8�͍�ڰJT�,�N ("��~��k�2C�6���Oϱ�q2X� SZ�)LD��*ʵ�6�7���b��F%9��I�N�B�u{�ȶ�{1���9TIB�Aw/��3h����뒧Lm<�@��q[0�U2a�lB��4����"� ���*�3�Q½%�5���;��{v 騴� ��F�W�/� �N��i�'^ʸH��ϵc����s!>�#�SKE�c�p9IR����	�ȫY.s�$��y,�k���č�b��t�B�V6�h�e+f����d_P����]��䨊�|k�ۃ��1#!N�gAN2z���2p�ِ���:���Fk�sU6T?����c�� ���W+�S�����m�9����D�.�x ��V��?:{�+�`���OgĬ����Z7��'�ݫ%g��Z�oz! �,���]o� ��}#S�{+1X�;q�����DFQ�ZC�S�Gx�װQ�Zd;���B7h�q��{�#����C��j�����^�i���6.jh��]��g�l���/ê�l�{��(�1�V"�:��〃��H��w$:�ܧY��[�&�u+e�ɘ�K�N�yx^��U�ߺ ��{�
�<'Um;> ������c)��֠B2���4X����8�e�3EC|���	��kL��}h�g��
8�P�%%��XDwd�r�m�֩ew�� ߴ�86���2���c�����^��D�6�ůyR�O��K�׭��\��;�	~sߙ�����+�"t�-R� ��Uw4U�W��v��.D��ph���&��3�6���|n1�ęzȫŀ��ۉ���~QU$3Fň2��S��W����~�h�\�_'j)T�Q�'��&=��難+����kS�*��[<����Y�
�R=�������-ᣛ����Ξ���X��g��A�<R\���'J���Pbέ��N��ȑ:o��xj	R��'>g�QS@AN�_ֳ�%���T3^G�g���wz"��|/��f~nֈ+�#�F��BT9F�w�.D�~�@~
���L}�v<��lI-��ž���GV�ۗRU�CR7
�'�λ�1�;�1)��yJ3Q���fL��8���:�dzH
?���*ey����U�/$H�������$H�@w��eg�ק��B�4h�Q��ѹ��0Y^��(�����t��nn�$Eū?���u��4m�i��y5*åژ9 L��E��@�ppѺh�E�d�@��c��hO�>�|"�h0����D���mT �7u}��D�����V�����s�*}�yh2�N='j�Stj�9ܿwZ��b���8j�����BN��Ԅ\9Z�c�r\�׫#M�Í�U���ڒ�0��)�`B�$B�'�n�L�eV�r�>��=�p�1�e&5���.��$�'�;�	Vt>�Y	.��F÷0�g�~��1'k�����Jɍr,��{{���o�a�_�Z?M����Oa�lt���h�[0�(�G!��z�c�1T�&~�k���+�l��Y�p�+�]�a�\ֱ>���*�uEz��/��Y��	11�~O����PF�s��bi���5�4�{Y�BCN3��4l�:��S"n���"=����	s�0��P���7�t��M70ZK�7b���ȭ1�6~F���D��uB�S��`��<$b�![��� c��`����B���v�N�(�ewl� �1�w��8��2\�\C\a�P�0�k?�8&:�D��d9�D�W0���G!�� 	]�ڼM�V��P)�X���������)K��#�D�U��S���f/1Li@�8d~�5.O\����M����|�|�M����t`nɋ��x����Ŗ�PYW����Ş���m<�2���F܅t:99��~��\�cF_��p�m�j��m���ܘ'4�q�����ܐM��"�3�L?�Hp_�oĹ�c������X����	,��3�5�zJ4��M�ַf��K��H}	V}�&�ٓ6}\�$���ׅ��L�D�'L|�Th�oS�T��C`3�;Uw�/��������!kcR�"81J.<]cw�@Wt_�L�A��1Bvlӻ]��Y^�������W�rd�hu��=ꛃ���4?�*i.B�A+n/A8�J/��0׾�.����)����1,K-S���i ��	���4��)8�Q�[XN�����ﰬLK���*�p�l��i����B H��h�leo�oU*,�g�#��=ZYF�cr�|�*H�~;��kά"*�f�$b���������Q�>�N���4��l�`<鄖d��% �e-���2gڨ�8l�}FfnjX���<��j�Ⱥn9�zQb�An�g��r�M�,��;r�X4�)���b��<A��w��o��nk����E˲�#���0�(��xѷ�Q��_xh�\�l��!��,Qa*�����F��Z%!��W5R��*r_��L!B\�W���h�y���
>�RI��,/u1�5Tt�i��tV�r+6���;0d���E�x;&u����=R�*ޛՒ�w���	]ؔ|˜�Y�ꕶ���@_5zB�1k)�}�0���J���3�	�ң¯dk�\��޾V#��UՎ��_�����hr���z
����_Z;�ބ����pl+�t�c5��׀i	��mvG3�){D�y�!
�GW��,��-Y�GDZ@MP��W� ��kZt�N�@ۯc�����Ҁs{ckbH�5PYi�@!J.y��8�N����3�<�^(z��ҴZ(��_14��X�e�7=)]�����ɏ^p�AX��C	\÷�
3Jf�KȌ������c��CJ�w�R�������t��v��;@u�R�ě�(<Ӊ��652UC�#��w��h��s9��2�Ѕy�	��X���.b��5�Q���/�H��L� 2�)+�f���:�eG
���0��-���b|p���|! �%��V0G�#���$N׵g�3�N��:�S���	���z�̇階�/�̹�
�wh=�W=�X1����!�j�O�Yh,�{���^=ySջq��ni��1����Α�t� a�%`�@o;x��ݐ2�sS	��K7�s	0n^�'",0���ͬ@(�ym? �;	�<�'j���H�u5��>����lC./W�B��r�'G��6n>#O���!��Ciߍ ���=�u8��g�9�c�e�=S�ˀ�'OWd3���l�� N�BQF��S��vZ��_�Up°!V���`� ���[Ā�w��(��"|ݜ0��j]�g'l��+����w��.�bՌ�-��"H+�-:�$8v1�WP̙�k�Wy3u��&f�7m)� ����>@���S���tq�ڙ�m�����@-�����G��f5؝o�3�Ԗ(JL�O�ɒ�tݴ���#���O\��bwQ�[��*��֜�E�!��ԗ{a�8p�a\D.��[3���,����oj��{������`�bF�q���}X��gQ��2��d_kKbo��f��0#��La��h$�vB�r��^���AG�BO�=�q-?�2֥�њ����&�Ȕ`=�A���N.�N��+%Dg�0U���NBg�,��|Vd->�\EC��5���	�D
�_�n�)@��9�]@�Z ����^�1�l�#49��@��.��mYrj��]�pH�.o��w���4$8�T�Y	���@*)U��w���X"�¶Qi��u��G��C^�jj0�=3��Z��әe��nl���3��rP���co��Q��!���[/�|Q���zҧ��X��.N�����L�VMBؼy�#��Tc/z�D�ח���AUv]�H�ev�g��-�'Ҿ �i&��Ñ�F�=���CȔ��Ɋ��m@����>����D2[�gʜL73ah}�0��u��o��Mc�4��òˋ��9�aztZxG�3n�ahnLh�G��O4�uH �^��<�A7�AvK܇du�D83z���N�����NkL:n�W�!(�u���p⇹N���(�wR��I���Ȍ�H�0L8�Z������,e��s��J�-,�*N��\4m��hG��r�5eE2�t�UR��3�5՝A�۠^����b�z5^~�=����[�|�y���p���m�Q��/}�����G�+�~������$�$\)���|�(l o�p`�Op�^��A��zƙ9�7[�>���b��0�{�S�y\83�u*�AB�Wi�=
$����x�s�}ƪ̺���礓�#zU����/F�++��5�x�<�獜#�r��\��<j@J3~�
C�mѣ�[Z�c�JJr���G���D��׹����IsC=�p�$��"w�f6o��ެ�rD��֙�e��qPv��	M����):Pz���y�`��J�ƅ�V'��{��J�JD@�|�.�����ۃ@ǋf��}�	 �+f^�!�������"X:`�iL���9��o��;=�۸���ȅf�N4���(hҘ}�-���"�َ�(��ވ_sV���wAZ����*gǨ{aKZ��ݴ��3Y|#�y�5���{;��\�_����SEYO�������-nC�b�hԉ@6X�D܄
�>�!��������}lroV�2H��a�Db#�V��F8X�p ��7Ȏy6��]���Ѷ[�uS�c���w�ꀑ�[��Z�c��=I�"uB^4�ցM�%��vӺ�\-q!6������n��u����eq��Z�3N2�mK�ɠ���I��	_��*[RHl��g��"u߸��6l2��&&pX�Vf�'QA}'p�8���S�?I,/!��G$�s�U@:w���T�&o�ӄ/�'�n�H��F��:yV-���I�SQx�0��ZK�܅b�t��,���f'F�<����^����n2^AK4��/���R`�[|�l��<�cn�Ir#���]B��1�%?y�p�O\���w��V,��PUYx*�
.�x
�>�}��ٛ��n���_0>�A��<�ā�U��H$v����n�Y�_�ھg��:E>c7�r)�m��$HXs�=���xj�g�dQGa��؀�M$�[��{��v�y}�������%�)2oi���@ٱ;�M���tHK�6i�ybfN���~x��6,�JUzo)�AB����!�p�%�����Ei�&��(��>͉��/�@��k�����.gn��/x}ZS̅�F�vG�O�c�x|�g�DB(��Λx;f��U�iF��X�J��P\a]J�Ӏ�0�8�����,bR���^ȉz� ��0C�Dh�����3g��$�@�m�`r�"��XZM�%�y�TX�6���G�d�ZEs�,ܵ�9'!!���s�j�aP�~LHB�u��s@�æ����j���sFg4�� ��d��OM�����."�M�s��"�e� �4hCdͻ ��� �:6�$����z�����M�Y�EmP'�V�e��A�ʮU��I��������|@���e�/�M� R���t��X��N�]-9����I&�|�N4,}��$��倚�+�.}���{c0#�u��l�{�}@
����X^3S|x�'���jI��ԹOD<[��n���7�O�t�'O�/8��H5��4r��fcpI�OG��Z�Q6
�4�h�lӕB����%?u@�T(s����<�i��J�x�gЀD���UX=3��1��.��ˁ([�q��$��;��9�2��cm
����n�w����n���&R����>W�d�|��C��mՃ�<���,�|�DN.-�Z�i���eNƴ4s�zvP��TI`=������x�^���.�θ�4 �_՚^�U#���;L�,Ԁ@�d�j�g=%�g��]�2ZJDM o7��T���0���r�'{�s@
�TYk�@M�ḛLx���f��G[�"�h��t�����ǉ��>�1�'M��<���W^,������GM?��_�G)=Zh7~����jd�[9�6�2����2��:�DL���o�}<��l�H�<�[�2��|L.�LW)@�Q7U(\�w�(�j����Q>?����U
<γ��8%w42F9ֲ��zւׄ���r_|M��}B_�IK>д|B!N@;�r�����VaZ_l-2xؗ�No%,b	���N�&0����j���~n�p�Y�}=L�n��b��6n���	�s��[�T�V�;>�'�u�z�5��-A�@��f-��`0�a�=N5�g�R���g�����3>,�QUAm�Fhn���$�����+�6H���2n���k�w�|�7B�ω�Ve��Q��C�LY6�Ȣ��O���ȑ�w�b�I�*[�i%g<Mh(l�)������a�r��	�k���?�QXğ�c��a��&�L9�<g�T�%�f�To��ut!���a��Eb����1�XH���$��5��5�R����|=Jz���I�isJm���Oz�`p�ñ뎍�>�{vU��Tx�Ё=d�X#daAx��B[T�N��;��F�G�9\��5�X$cNOz��[������pR1� �~�5)���/�J~����zWxC���b4X�p�6Bz�GtxM������(L�ô��Ž�����j��k*��!L=���[�*�Ǝ�o��%3���ӑ
��{4t'�f'�J�r������0'K�T_�L&��6}���D#xmQ�~B�����B�(+@�_L1�
��D����^g�(�.k �i��Ȓό�,�u��c�	�*9���o�]�깞�&�
��?�B��	mtA9�E����q�Y��G�D�e�:m(��a�R���7>����g����x\��Ʊ�>-��[�M�9�.T�`�d�lt�$L���\Uc��y��m���O4�̃��H�d��� {��� �=Q�K�i�h���&�rB���@l%ӲS[�a�~Of�`��vW݉Bto_��To I�����{���؀��sW���=��&��@�vO�07x��ϸ�O�=D�v.�Ѿ�|��㍃9�q�����FsJ;U-�ςb��}��|Ys���(���@̅+=/���A���F�"�L�b�8���h,V_j�e����0���`u���qucj�Q�����i(����G���b ' K��Z��gch�SVq�y1�v�4J��!1���=v�k�^�+h�H��yt���H�&��M��U4i��Ѿ��d�U���G��sԒ�ػ�iF��=�Y [�zn�ђ���{<����զ��P�=5v����yT�7_���<o�=TN���)2���`œ+�l���Z�寞qo��nh�C���*ed>��p�d˫9G9����m(aFӻ�O���G�C����*��oM�h�+��?��}��É���b������F��@���B�������8���Y��"v=�h�:QzL$��ɫr�����0҂=���ѬI��x�_-�X�	�i[w�vtX���,}����S#�)�|��b��{�d�xϛ��0[�TU�,������[�n�7�_�v�
��_�K�`c�)��a��AH����s�'ʑr�
s�*oN1�$m?��/��(Z���S�&H�֤�$Q��@�^�,ʲ�������4�;��f��٫~��u��܍U{�+���������{�q�oՙ�5�ȹ�k�{��>ē���Iu�$�^��I���-h� zt:֘͠�P�� 7��<�X~ŬF	h�:Y!�]��`�Q�@��J4oY���]��)7���v��`R�a+���x���{�|�^��1.�j�N�v��pMo�L��ۣ�����K?Xc�xZm� Ff��Hj�IG���z��sl�Q���}�}��ѳ��l8�
��JM�rڒP�/�}5/�\H3��]������"��A��_t�dsI?�m���{�2������ �`�e��ďF��IHeT1��eP���Q�[Q�p=dN�R z��6m���|����n��p'��S���o9oZ"b&����G|#=Mn4��m+6C9H�W`u>�?찕Cūa�u^VM����c��|�p���X7�B�8��m�/L$w]�S7?�8���m��$��9�g�$�OQ�f�P��^ç��0��+�C��U�U�L�x�,�A��V#.-m��#�9�Na�Ea��5��:ӓ�j����˦28[��I�"�~w6��c���=.�}�d�s��G�:H>ƕ�f���
8qq�/jɞ�J��Hu]5��Ĵ2( �͢._[k�;�*��74=Y�hn����bq��pH�&šKn�s.Q`Zxe�)��)r���?��CX׉�?V��&�պ�X�����V��r �}���Z��V1�O�(���8"iY$���	-j��,�Ɓ�<P7��FW�0'V\
�5[E��H4'm�I���B�XL~mX�W�BT'�|��)��F!P��A;���:��d��P`�]���z�,���o��vy��)RuJ�	X�+�"�
���x;���]���c�����r����G9ȋ�zSH;	���%�cv�@C}W��IZ��1��Dt��2���ߢѫ�zOOQr�*욨!u�`�t>n����$��hc��_:x���s[cjF�,R)�`� ڰy�aK0I.:�H��,���`�R�+�k��������v��`��pX���;�܇��[T�����D��)Q�����A��8| �^��6[�R�,y���� ��h���*v9���VӾ�s���?)�B��j_��z�T�i�&��Z7�f��d;�,��yU��Q�1P�I@�$sc|��_Z����p�Hʴ�/����s!1��Y������h��z ��ER����w�^�1�Ƙ�Q���N�-��\���{�V��_tL����Z���t )�����6HR�P�96��"+�^[���=]�n��Z&	K�L�����ǅ�sG�u��z��v��w�Σ|��R�,��m�1���z-X�1��ފ�gk\{ޣ^}R|q�(1�S�ED�a�Nt�$
�N����S���t�q9��l��Ph��r���K�]	�,����N�>�s1 �m��->��G�O���c�����M��E�6�6*�#^E��Ԧ���'u��L�>�Z�E�s؉8��|g�� ��i Un�$,azw-�*�9�/�7�c֠�ʒ�b�oI�m�wJ�A# �4�넪^�&ۄ�#v#o�?v��s�b��O%���珦��ȁڥ�n�����PL���������ޠ^��S�-�In��>+7���cjr~�*F0�+�AՃY��b�(�ְ���p�N��-�@��[��,z����̗_�[M#+�k�yuD�lE�(��
b철�
)'�D$:{�&��o��k"8L~|�(:��|D�����347PT�+¬�\9!��aA �\>w܅����IB�z��U1o�V�TP5���<~�v��Τ��%��U�O�	��rS�Q�w��o��6�n`"��n8PJȞ���iYo9�1Vg�:IK�޶�8��ڮ.���P�7���^�51�F��ט^
�����q�i���� ����h_C���C(�&W�F2\�oe���&z�B�Ԙ��$�l�R˿B��99o�#I����S����26�"�����e�]��{��;<;�y�.�n�	����1.3��ڪ�n�*0m�If���T��h�G	���S=R���o4*��-
ϫ���B�-�D�O!�����q.�MC`���afZ�Ճ�Z�W�-x�8��&�S���������N�$�{�˜2�j?C'��b�x��D\��/B�6��tk׬!ǏpK3u�N��A�[�R�Ċ�ZL"����Ż�����S=H��e��ݸ��
j�ie)t��z�'.����{,@�E���)����F��F���U�* �x�5Œ�
����]��=�Ql�0�j�.P�V���4k��C�l��x�u5df�2�a�t�\H)��Ws�6x�w����B��@4^���1��?���2*��A\�\�9�Ϥ1T	�4M�z<mɩC�<�U:�e�[7r�M�S�u��}s�����Њ�*)�����n�}��KxF.�(_7��Ļ�����J�0��O���$p��j3O�0��ӄn[,2�q�7��ْQPm�����P�<Zþ����o�ܦ^u�����ȄV/����{��.k�u���M� �h�{Mb�A!�,{����	Z^��p�/���G�V#��*��]�rʡ�ft-��oa{���Fq��O�l��̀��&ۜq'��)���y�9��~���3�o.�:ӹ���kb$���Թ�4u�y3{�[t��c������s��t���#����xe�p��տ��a2{0��j`a~��Pgt3�NO�����t��At��L�􆭠���`���Nw�J���y�>�	6$3꯸}f���2�ab"J#-%�zN�SW�ÿLM�Z����J׻*�B39��>�ԫyR�1�AD��E`͸̑��cW�Y�U`cI�{5�܊�큜|����_�M̆0f�p��غ��M'T?�S�g�0b��n�Eg;�Ո�m/�O�(n#��s��7A\ɹ��T�� ~QK��a\���+�Di��o�B�'��D�^ALM$*Z��D�-f���y����(��ҡ,��K[�ǐ��;���Ȱ�.��Ø��5����,bE$U�瀞]e��p����~OUp�[�*+�.w��z�3�gr���n�!wV����X�U�Y��M�5j��%��|����-.x�:o}�������AW�qy0�b�nI�Y�SL�����!�v�"��]-��~�+��9��Ls���z��5K �\�B>Bk~�y7�RL�!�1��{qY�CF�Ӭ��`�Pۍt�O5�9&~��v{�B�Ey���hL��K&���D�q[@}���4+��N�**X�e�g�Ң��Gd��C��a�%��(bsvD�����G�}�	0%���Ӡ��*�USڐ���l�"��$�ۑ����zYr��~fā6�D�W���:��H����';�@_�*�Q&Ň�q�W���bV�P��[X���%k�o^��wr1��^D��^�W��r��G�~K��ʫ@j�t@����jF�3:i}��k[6~��A�zŉ���
�/��#T࡮��`�o�'"7�"鷿��tXmVvy�z宰�	hAQdH�-1~z�(imFD����c�8yQ۪b�� N�1Ɯ|��?����:� �!�@��TP�g�S$~�w�k}�Cdn$�MIŘJ�¿]��bH�+��Q��Nn�w�Ec�|s�]X�ߗ6��T6Wç�O�ɝ �	�u�D��:�Z��lS���XEˇҪ�K(O�/�٪�����
�e"�c�"�~�t�cl1�������kŽ�7#%F�埓���6IJ"�y{����5�V���Á�&�hԧl�v�qq����gi�7Kf��$�u�u\ [b�����n˃�3B��N��ʾ�͂�S'���	����!�آ3�C�\�z��*W�9g�q}I��Vp
0���ovg���Z�w�D�k���Q�]�+���//�g���H��c�h���Z|pǸ��E��|��rI�����8���4��$��֤�{�����(��M����k*�v��'�!N/�{'Q���ѓ�z��n{t��a�ѫ����7>�*�x5�h}LKY酤~c�>�ϛ+�<�kF,f��`Q�@b*z���5�W�U)8�������+&�7�l��G�K. ��x�qhD���ȃ��#A�Bbv��;�5��flH��:���1װw$HM#@@� N�a�:Z�%<ߖ�Z���Fdl�]$�=C�z�Hp~>t��f��P{i�Ƙ�� эE�_b7�y��9rz��L�u$in���*���Й�7�6��/=���|;�1�����埚Bs�5����`D��h~eh^�k1V]�8+m���6�'�\E��6�I-�����L:��}�ԃҷ�VGWƥ5I�����<�b��v8�܅T�{)S��=/:�=�>�,���f��~p�bR���p�_�Pr/�Wh��Pٳؠ��[6lK�Jp�R<
n@UT���iۃ��V���X��RQ�K��2����]��tג](�C���p���U�wP��<Z������D{�U�-������R�q��]�؏,4���@)/ꭓ�q���/��$��Lƫj�d���ٞ��� Zm� @Fۿi:l�5�[��""ޡM_�J���=��n*Y;�/�m�����:�U����J�3�h��_(C4�7��=�n9YD�9.�:֫���K	y��bS_D�j{�"?Ώ$x�����p���?��e
���(y�`|���@~�_��`��L�	X�ٻ27)��_ �������4@�!!I���CV��r���˳�Һʻ��r.f�]ߨ����Qn5\�X���ҀAND��+����y��,���2��a���~{�u���ّ
I9�]ϙ8��#Rom`��c���5�'or�jG��)�#�D��K�(�Ѓ<�� ��'?�x��aZ����,h{��b>�NV�F��m�ǲ�~�x�2�(�/����`�F�Kܲ�����\<q�������ѣ���P�� g��`��L����D�:8�����)�S��8GT��JHt��O�l�.�X�[/!��&�ЬH���rϡ�Ԕ�}L�L��5(^�-�v��_�)�ow�p��A�@���T����F�Y��Gy\OЈQ��P�;lv�L�k�a���$�<�� xϠ)Q�$���n�V���0��p�G�Z�p#��N�Ȋ��� �pWi��/�۔�Ȭ�����C�<�q�?�c�Mݒ�����#;Y�g�~�v)���$>Z+�x��7��W�ɯfx�G�`R lW�ڌD�1��&�]�r�L`����-\��G�Fx!�g���n�M���ѹ�U\�MG(ѡb2��J�7�-:JI3�������T�G�E�`T��-˼gd�������pachfŔ�w��
�N,gr��ҕTlh�����x��~���켩ƫ�#"�|��uπLؽ������?ZT�Z�A('m}Q4��w7ܾ���f�P��^��T+�1=�T�I�:�	˪�#��~<U����^�8-��q��!l5vtն����9.SM�7��M䱸떔��/U��<�����\��H��J'�x}��|�f�Z��S���$,��l4 _������5h��6���hg�to��؞1n����C�>^p�6M�"2]��� �!v3��(�y@2���^�9�h�����q�z�d2�|���E;����[N�=�����c�d�T���F�h\�3�������`P`�˳�K�£k�;!��<k0$�#�bQE*�)��:R�{/��I���7���6y����w4A;�m��Pt�1[�&��������N��.	�'/��an�Fp|���������j/��n�Y�f��@	>�uG_l��p����/��tH��AAh��%��E��GiEk�)�YdX����~�~nR[y�S�
��Q�-.q����=���/��P9�Yķ����)���Ѯ�}��~�>r�ف�5N����q��S����M`��`4�Ϧ�z+�S�Qe�
{�^6~�F1���ig}>W��m1Dm�uA�����������]1۟��$�D�ei�����H�ky�k/*���og/H�;�#(4^Ř����)Η���9��V�[";|T��2�%fC�t����߲Pg�NDK�Y�껌=�*@! ��H
(f�h;Δ �(d�b�0>��,K�,1SAD�|b]:;_{�U��o�"rcZs���Mz��b+3{q�Xu.�2�Ei]l4z ��C:j��ZM��U_�>_����פ����2��@#��8��_�r:�W{��S{	"�1~U J-ƈMIN�L?��s��.�xGkKէ@�go~��F`�YB2�Jw��C~v C���܁2�"ǰ6G.� �����e!����7q��X��"I〥��(��!�|05�AS �[)��u��l;N#;
U+ss����0��U��t�Ҋ�n.�浇o�m6 UL���Z��=e���[^����"l�� ��g���b5�ğ����Xes؄,�]v�
��l������ �ٲ+Vpy�g�폶��D� ���~���^	�oF�Vo
�'�\��g�a�ʘټ�YDe���.��h�/�T�n��)�(0&ek�I����^T
����.,�z�_v�(���n鲁�MBA� Β.��� �:.(0�2�S��u�w;���֞�,[a]߈qj��Y�  �ZR G�K�'����5˲�Z���p�J���9P��?b�k\�l"'"r?�{��1Q��3
ܒ4�K�J�>�[b�������R�a�ڧ���nT�!��������z�YS%k1�V��� ���; �ҽ4�_�LqJ���F�#+^~
��X��r�Z�@ةИ� � xI��f ����M2��(c�Z��T���۸k]֞��`�Y��Q��>�!��K���^b��9U;h��%>�r�82����(�.-pSxs��c��Ԣ��!]f���tt4���ra����:�U4���^&�����!ؿ�$��t>Jz��+ů<!"�n�<�5Mm�;�Y��C:ǀ�/����3����n��X��W����!޵��H<PN�f�G�.<�J��J>x	�;�{�sz�$�d+���4��K�%<R^{�`H�1J'� e��{��^&��٬�Џ=��a�i#FiGBu����3�%�4��G�Cl]�.��ir$]'a�W�b ����,�h3���)�߱��$-c��[B�x���j�z�)���9�Ɏ� $`a�Zq���|ܕ�ST^�i�dOl�*�Ȇ\J�8���.��"����Vk��&7�"A�};����߈R�V@�l}��	��i�y{g./��2��g��h�d3D8�Ԙ7r���&�HlZwfVB���8쁴C�=p�z��*߇��Qoc���N�mӜ�1��9(Ο���+6�V�	r;~)�F;��v϶��&�0�y�(E�� ��nn2wr'��j���aR�=�M����B߄��@ӆ�Il�9K�(�����vL��WԷg�	���jU��X�H[�9إrwn�F_C-�a/VJ>ZR%L������Վ�[p&�<��VFǕ:����^��C��n�a����Dr}y���ړy��Hj��?�����Nu���'��ȹ�w��҈b�˾��{�uWN��]x�EA�J�h.�������l^L��J��y:�H�����T���n�髠W��������sí��n�u�m�F��ǅ��#us~;��"`�ҭ�)XV�V�L�^ՎV�sL)#�=��w��y�{��+�~�穲ԏ	�5��UaQ]�XV�݉*�m�\v,���St?��ז�%7*��y�P����O�S�?oF��18�^(�@��a{�WkrQ�ŏ�I�<uE>��� ږwSM?Y��M��^N�2ᵣ��2���4I�;}esy���0,����vb�8@���~8�q�i�^� �Ӫ��a��mЏ�Km���2�'��H�PN��(�DF
ԧ����G�,�P{�k���b�� �#���)b�G����ő(2��ym����^i*5�G�%�p��uQ��2�Ւ���{�8q(�鑣Ns<S�����R���V�G�q�1h�Α�x���7Y���9�������ѳ��\�<�ǮF{��Lݯ�em�#}����P���(�l��bu�w�kj��Bj�{��b>������f�<:�j�g~w�"L�c��k���0�>.�V|�����Ӯ�E�Øp�8|�5��n.���#���e�=ݧ&\�HLrK3�usHa����o�*��[��,�A0L �y"~�i�=b�.�/}����E�8�ճai����W��'�Lr|ޞ|��;-�GV׀o�"���	~u�J˨�ؑ�f;�Id�g���̝�PN�n>}ᕵ��?Z3��ϗ�fnM�Fp0�4m�ON+@
�?��>�j�m��T뚙�z@�7�����cXƒf���5A�N}>�0G�;a��:��{+G ���x�Fi �W%m%���l᜾j�ܭ�Q~hO �W��u�s��6t� �]�����4��+�ș^A辩 ����ԶV��#r�Yl�*;f�j�y_p�Ǧ�*�d�Пt.s��]+��V�!Q�5m���.%H>�j�+��8�!���xW��J����ꤰC��t"�񝰅&d�S���i�$�'���a����|I��*|l�XGG�E&��t�ۄ����Q2l��NǶq,�i�i;>�1����ǜ�P �oW>��q��Cٟ��lD��A��6�W�F�q�=��h6�o��I^3��M+*[���Εײvt\�(�gؒ�	�2Z+�����\!KG>���t���-\pJ�S�`�AZ��ҝ��#ׇ��1�(��[�f��1ch}�K���a����x@��^�k�%��Qx�y�G�տ|��Ip�}�~8�x�s$�u�j�Yʲ�R���}�9�8���1l.7�L&��"������DB��=	��Ƀ�	p>Q��g	Du�3���]=��j=�Z3�aŔ�W���A{���)�#U�\o�> 	��6]��i���_:g7R�Z0�+����*D��u�dy���c{��We!�T�h����V�T���N��5��2�+���^�=i�`��]A)߭LL�i4��w�
��Aoֈ@
��| ���K�Zb��W�S�������h�mu�G�{�ԸI�{IQ	��㪪`��j��Dehj|�>�`��`�`b�	 ���>"�©,�*�ex���Y3tSZ]]�����f����1j�̱��n{�{���(�h�,ظ�����v ks��"܁�
��!�aU�X�Z=�hw��y{�_���UM~�o�㖉e$%*O�[S&�%ݦ/���u�8VyH �QՁ�N��d��
����-��;�mE|���9����=(D�g�n��®�ii�_��&MJ�ڬ��\u-��pNF�J�k�,
Д@4Wt��k H[�����p�Y~R��}�M��d4�ݺ��Q{˩'���X�K�(�p�C\Z˪�T��7�*��[��Bٚ5��5
GqZ�6���K�l�H%n�z��\}$2!+� �w���=I)j���#GFL*���j�I��P�[=��^���=DW6~E��u����2��nh)��+���d�;;�_�ރ-���`@��'�>ň
J����Pu�3�X�H�%;����� �����vZξ&h�S�7(�$��>�i�����������6��Ju6�3Khx�U��K�c+EIi�L/I��L���5��@��PEE�Ȫ3�Ľ�B����>Β���z\�O�@�m,o�IMқG�]�/�G�^��{.�49=haɠ\5n�8L�t�"��B��D*>R�k.#�d��ڊk����B��`�v�A{�DUŝ���E҂��`�����F�Q|���2T{	���`DDfV�dS$5	���#�o��5�r(�������������{q��-��I�|�#�'�sKf&�}��	�d3�3��*��:����!&>~��w����i}�5�1C|�!�?CG��1!S��O)��Wi�̃�x\�*�޶(�"/4K�f~<�rO���K�t�r�R�Tlx�����|�d���y_�;} 	$=��ƒ��_MI���/�F䊇ؙ�˷�1�/��#Vz�V #����m7�+�3HW�ɡj�ĞE�)�6����~�����Q	;�|/���o`�;�80�9`<"%$A��f�ߩj�M;�G,�[=�[���E�9/������w��A�вx��	��<�j��d���SK�\\�)�nHl����(_̾|K�U}gM"Ղ�)��b
��2Q`�I+<����߭�S�Z��<MJl��q� ��ep��)m_����f�r������CU!)%�6��=D50�\��M��G�pݎ]�Nl�	o�n���Q���`t�>�F.;\B��i-J뗮���j�2�c!�n�V����ml�Er�[BJ����DKt;Y��ߴҰ��#2'�l�2��M���"��	z6�mt�S�9��r%ov�<WX3�vj)�����b�ޝ6�I�G.����w�.�c��9i>�#O�C�⋛�˸�� m��|�:GR�ُw�{3��(H���Fw�������_J��3 �w��ǁc�%-OWF�,̰7rڷ!쥧'U�e�5�iGy=��T������T2�B�ز���0<���O �|/HP|��,x���
lA��|!��'��n��O��*^j�
q��ިO��+ȁ��L؁�����k�K��t��K-e|��:囔�#��)/��������Zd��q�*�����E�ꨣO����$3�(17K��۰�CBQG�>$��
�@� �fm<V����2@�U"����Bs���jݟ�di��Hs�}2��6������$��Y|�j@� ?=r�T<�P}h@6+�M�2�+w�m%�#��ӎ��Tcs=8��+f� g/\e�����ŉ�N K�<�� ?V
�/Q�s>�[�ۡ����&3�#N�|����d]oMES�@dz�zvC�ˊ:[ww�k��FFSCȬ�[琹� 6�u�L�;ڜN����?n5,o��c�D�\|Κ�j�t"�"k�������Kj����;�)6a����-�7��6�'ȣ�*ԗp����I��/[T�?r��1�f�^�B�PB�Ŵ���-���	�=Rr�#�ؐ������܀+e�}Kk��������i�	������{�����!Z�{l��T�D$�r��9�I�>�sg	���3Wn���K� .h�����SA�P�ϐ����J=. �f�r�ʮ�P	�w�?G?��E�K�DpT[�y/"K�D�Z��>��ȣ�T��)T�C���6����..�øŞ��['����^���u}@�.J�Q���v�pU�4�{X�;F��Ic�"���Y���{F(]���V)(���C�ȏŁf�� aZ(�"�3_�s���`R8�$ζ�\j���/��x�Oj �/X�������*F *����ZU4��2�޼��nt���ͯ%iB�)z徒�o�I�4�ocM�w��`��^V��_:��N,���moHz�B�')���C�C���}�9�����6�t^ ue��}���b���Z$�@ǰ�����db
*2��M�vlr^�&/V�y��4� F�$�&���1�ȡ>S���{՞^���cM�a�����w[���]�p7H3u���yqXb��������_q� �.ҘD��C5���r�%�۴"j���X!�݂�6��/;xi?�8QaX����q��l��d�ҳ�Sg�� �}�|�
n8k/��>��|�߉$}`n���V�ze5�dW�{�4=��T�֜dB�`�أ"&��Q��W�,;5�&@jk�.����f	f~�^:�M�:�a�.J�;�w}9?e�Q�w<M���:���@e�F�s����xK�<����Vp���N��i���]�,��Z����N��
=��_�>TM�(����S4��15z��54�m�J�� �~���Fr��lʾ�H�â��5�Ю�ҝ\�E.��h�c�/C�JW��U��w�1�,�G'9�������\�Q�MH�YA �i�+<k#=t�2�7�����H�I+�Ks	Ad^8u78>a``-"%��k�����}
�ؒD���t���	�ɢ���s�H_zn[�qo���R����8�U-���vtiW1�Tr�3��`���kf��λ*�l��q��R$?kmQ���tT^�NF�wb)�i����+2�^VI�~Y��t.���5���q�R�Ȉ���s]�A��I��,�q4�]W��^�'X$)Bq@���no#'���⡳Mg�`X��|MΡ��������%	�|L��Œ,�i`��+�d��Y����1K����xW�u�"7�c�#�xܕ,���W@�1�܁��aL�Nc�R)��� ��,2,��]��f�,兿�]�UY͗2���D�l�庇��-B�&��]���|�Q�?��:��)��ŕjec~�BZ��q����.f����.�}\��	�_0� ��퐽n����x��������?��
�iE�$1� !�@�GUvSa��V��%���(C�>X�?aڹ�����2.��n�FU���K0ȥ����;�����m�}M}���Vg��:�w�r������U	��Ȣ���D(2�������~,�3���gs�e*߳;���Y��
���`��\�D�v�oY�E��J�d�BeØ0��1п��X(wSo+K�RIQGSJ�1MI�^E7`���M.���ñP�,H��{��*֍4�3��Ϣ���ñ�DK����~�*Lc��z�?�lt�3���]�D�f��?-�!�v�B\L7\��T�u��(�fm�!�t���&�����Ό^�9���?NV���k�~Ɗ:ʌ�8��ia TB8�7~�rń�9] X�/���x�`����Bb^�L7*��3��4�5��_E����ei�oy �>
�
��eӳ��Z~�W��=��4�\�`�4���j4��A����mlt�-��@��b�((I�ou�
�K�[���:p*�&1��&j
p�ω�!r�V��n���*�G[�s��S����<,�0֒x8릟�DD��`�O�Ij޲Z�O)7~�ʧ	�C��{4=�)�]%�.�B�ek'�Љ_C�ۉ�Z�%����ֹ�Y�	4ݿ��@�^vlc����xh�j�Bxk�^0��j1��y�xO�
|�|3�� ��1k렷�g�5�\6.TB6��|���ဲ�[R�$KJ�t��\,f�������J�"1ĉ5�9F��D+����D�T>DшU.M�ُA�	�ϱ��,un>�.Ɉ7RM*e�`P�|.+*���;�]I���v��r��Z�W�#��Hz\������po���� �|Rm��Tر�#��~O#���[�])�?�@馯���59J8!�`��$�+h#��8�f�"X��x�ku9Z��8}:���ć;:�E����R���Ե~3�&��
�O?��������Sފ"��$���[H�
ġP�����$r�k�t�Of߆ۻk�?6�����l�q�&�Y2^<~��`>�Ȅ��-2��	D��W�x��mW��rb�y���H"�P�g�f���U�Z/ڟKT�J}k�b���!���+�R��� ^߈����ͨꛪ&�,�eI�Q�P%Y[��Z�#<�~T11f3U���C�jX�>&�W�2���?��YN��_5��
~������ʲ�#Li�4���9�x���ڽ�8���Y�ē���	�0~Y�lݫ
c�i�j#���s�2�E^��D�o��~cf]���^��R��\�L�+Ic�D�辍n�a�"滋Sǁ����C:̢1����� ��07��&�E -~�i7��w��d:��T�W!R���b�&�!��Ji�!x�#������q���u�~�S�4�m���z��w��{bYީµ���֢��2��@?j&�E1����!����Ȕ�\���$��W�D+8��L�1����z�lI��V7AJ�@Z5�큜UQz�f"`&���q�.tjz��?N!b����枆yupJMf
�5�t;"WҬ���ƾX����+w��oG��*��'�Jl�O���XT��U��ya�TX�0�+M}���(�e��f3ݮ�xb�=:�7,���Z�^!t��-}�R�C���m�)�����cߥ,>a4o�6�F,=�$�y4C	_�H����Q��
5$�Z�*^]0,��-�Bj\J�"�oT�#�A�w�L�f,�Ktl��>��#e6���MI
�yRw9��A����݄�R)ă���(�^��|f�Mb{��/*�F�6Yw���� ��kǗ��㋯ʬ��k���fαs�;K�\�ׇA*E�d{lm�16�X�g~9����C���D���ל���.�Hi�k?���In>W��G^� ����^��^Ƴ��iD2I1]-cÔ(E_�v�X�֪>]D�HC2��x�K�h���s���ߣ����������<�h�Ot�oO�a��ӱr�Й������Z�$�<�.�ߗ��&�r���5؈�s��?t�@FQ-����#��/��/
ڑ���ק�'�[��g��_�a2(\�w��o�h�ƛ���e06�1������I�֯9�߫ryo*\�@}�n�UN���d�=7��'�fwu!�4K=��	Q��~���l���4g����N:�������i�L�ݱB�h�s�,����̫��ʊ����+d�+���C��ĕ����/(��p,��F�q����o��UX��rz��-�#,<ס�R5�$an�X�z��y�C�i�J�����*`��@J��p�Cρ��59�fmw��Ik&��W�z�C#sќ*��!=�D������;�I�����T5����Q��5٩������OJ�E��^���M�-Z>�q�ױڰ��,��"А�O�|E�y'��1���a��p�����D�7��Y�#��Y���T�����lc�@C�f���*F�V���2<j	$�%`Y�iUɯ���T���T�(�D��Å,Ά=��z�
u[6Y�k�=Y)q���`�P�O�yz~��'&��>����i��Ekό���n��,�۹���8���:S�Â
}Y�����~-�^ �{�v/��&;�` �1�84��cj�s4]U�߃q�^�E2����!��#�;V��~m�����8�4�I%�!K^᪒�e/fe�����& =�=X��/g���;8ɝyt4�� {&#	8��p,�3.�d�[��0A�z��#�p�U�?s�s6�7�9i<\P���l�T`W�{�_�\'�gO���:fk�������4�7:�<�~�^�C�S���U7cZ-"2�ܘQ�2nu2R����Lc@/B!3�Iu��-�TU�t�&s�M�݊$=�Q�	�j�LX���8R���X4����4��bc���K��cۦs��H7��Q���q��83�����E��G"o
K#�����GA�n#�y�z�/�W�{����u�e�>C`v��NbB��}7��<��������l��������"t>���!F��w��.僒*�V�^�F�����Hu���Fڱ�y}Г.�izFx���\�m�{o��&ܒ�� ����M�҇u$���D�l�ԸjRar��� ��p� v`�O1���§m��$�A�v�,L�-��fv�0	L�����S7�zq���Q�p�{5����l�4(����L��ҋ�%��h٩��.�8�֒�p����A����%8�r�U�˵���qM��M;V�N�{5�H��e\ZH�zw�l5��A�Q����a{Hx�q��:���V�ƺ1�q��Ω��'����ȸ'm��qZFǸ��$p&N2*Z#�ƭ��W����LԸ|'�/H�Q�r��H�J&ȧ��ZH�w`�ɾ��A�C�9ي�5j'����D�fX�\�}ڏ���qo�����V�=��A��~�3���������ȁx���&��8�*uMq���2�*�n=`��(�)�@�HI6����O���M�L=1�d���Ԣ���'$nv�?�Z�:_q�i�ըD�9]s���]�X�9��j�b�70� �{�}I�~�K6F�|y�f#N	�M�Lv.$Y�/V����R�7�����<(I3IIٺ���4m��~p�T��N>Q��~Zs����V����1��M�@�;���?BG�;P��}ۀ�b�׎�k7"��RH���֍4�="_�C?y�8�)���@ơ��ǯ	���6;i�m��$�XW~��j�*u$��w��o��s��[�ܐBH
�)��7%� 6��o���1��f�lڄ1����-�����T�(�Ȯ^>�o�ͿK�륍��5ʽ�*�� ��qI,c@�u; OL{��}M-��E�ރD|��$O:�{��)�|?�`e@�[U��aU��TȞ(ه�pH(=K �p�D����^�x�"��HD���j�V��:74��<�T��HXV���W�{�Q�`Yy}�	�4[���!?�ۣ�ET@$�5V���D:	XPs��"Pr��K�6��/@��@c��n�+������c#,\�z���[�?�h��T�tx��#}�|�[�a��^�K ������HrQ�}�
>�qG�½!З����沬'�wXIy�<����x5q�W#�����f5e������~q�(s��[(|��g�\ӐA��S�G�4E��s�۹`m{�aJk�2n|m��7Gd*�	��l��:A�R�$ a�"p��&��&E��"5�An���K��n ��2rx���C6ڞ�l>�%[����/��m�ʥäת<CV?�̤��m'�X	��5`��ԁ �U<0Ex�߸�l��jחZ7W���%ʏ�Ǿ���\�]�'#Ό�g��h�s��[0�e���1��+�6���������T������*8`�:��9��a_�,�!��*�τ�G��˩�>�A��p��� ��L�N�"�20�@�h=�N��)L��h���ݒ&��ի�>�ɣN�߮������J9Ț��$�M�.��>��ssP��������?n΢Tz�i;�ţ�M���}��z�?��J��u3�Oފ�@. ������x=�<b�|��5��q�P��A @����`��dJ������w>��H	�a�g��&M�n6�;��ә���Ƌd����P��'�֡v`�O�ηP��`6^�i�L�`�sz����<����S����<%}�WFbv�
��VT��~]���"�Dm7�DZ� �Z:"+�O���Mvz���=�w�1>I��� w� f�¼y��Aw��#�D�C�q�iit��v����,�O��B�����k���x��ꠄ3J���0u�{�_y�&Qo2W+!4T�S�_n�����tw�� YX]��78!N!K�g��C�LEg��E۸���!�����ڢ_��ߺ>6����)����22ZLA͢	W��C�����"2K�ձ�_��{�Y�`B1د{��a�D�<.0��B�<w�����ej�g�RsX�㻄Q�
�Z#�Nx���	a���kL��A�=�'2w����>�g%�WG�wp�R���M���c5��oK0Ƕ/�A�E����@�g����-�]��XBl��֡]�ڱ�����x�'c5ݠ���,�XօR}q�1p�@�?�'��yd��Ov�6�bQ\j\���p�A���*�+�G	�.�i����1���@Q�J��`\�{,�Do��>u�CL,}�VD��	-�m����<����O���ZIMT������ܙ�����¦�z�J>x,9�9g nK�V~�HM�-M|�O+e�Q]��;��6��,��3�&PpT��|<.+�xK¯%���"���^s"�2�W/�AxF�)�Oz�qIeS#0��rF$L�!��8�����ɿt�S��r���B�������W"*w3#AM ��mC�7�8��-r�a�?�&q(=��Ģv����{���{|o���B~��;�*HN��;ઈ|�K�S�U�Ϲ%)m�q�Mm.Ց��>������fZX�9t�=���J�Nxn�Hkap�!�9e/�*�,���D��f|���ڠ>�)�#�Q��n�<l�7%�Va�)�J�|4ʈ�7�i(r4�b�P���V%ӑ�t"(���� �rX����0����;��KU�K�����1$X�̼)Eī����ڡ��C�J�&h@3|N��$��L��*�r9�t�;�W���#�!9�"����4F��?�<617�nTE�=�u�	�3x��nI�Z:�&�.k�:
�����R��v�4�����#��v���6��t�[��r0��"ɀ�sf/�&\��0�^Ƙ��.�(�����MU,G��Z[���9LKH��``��Ey3gə^�v���]s�fuJ��舥��Un��W��Ϟ�kE\�#ks@
�R�	����<��k��|P�����"�HW�Jwo�|Ԩ�s���p�U6�m�G�Җ�:=`�n�u�+��;}���#M�=���1ڝ!��/�s�1����!�WF2����9=����?���6ժ/�١S1_H2�OsH\aO�`(d�4�����m�\�۵g}��'iÄ�40X��lD*k*4�c0?��V��4T�RǮ�!z��2���:��׆�'A)�C��g%f�V&-�5ĺǘǳ�e!�2�\��$T��PirU#/���_[ �8�S�˘?t�R���;c��P�.�O�FˡP�*(��Ÿ���Z��}���d�7�4Z��-&>9�$ �zV1GC'���"DP)z�W�:�����:!-��\���P�V�ԩ��z��$��\�O�"cf�c �l�S�n`��/�ʿib�P�؜*��V$����~^�[F�k���^���0=�2FR���]����r/��j�] ��]�>�8yp��;�Ɵ��SCz�j��ӳd��44ɪ�;����>]PnV���m����O�맯��($��fS�;y7Ͼh����lt�X[2��G���~
C�TE��\�Р���ƣ�zfuw�Bj���]�?.���k�Ҟ�?��U�h�h3�RG���m�ϐ�h{���'�k �ߩ�q�YU��u��W����
񔨄x�WK��u;��B�BtL�S��$�P|�?����&8�QOǳ�6����a��:w���'��I�.ȫ�f���w[��� s��k��*!4�h�p��&aj�r	dQ�&�����uD��5�?,	��� ��b*i9�(� ���t�ܮa��C��ej��*��/���[f�R���j�	�"�΢�����d���Tn+8}�H�T�,��A\U�ߖ��vF���TMl~��6�vO`���~C)�ߡ�ʭ6��W�ea�=���3mz{�!��,~��יYh�ͦh'��D��*������?����ay睳T�Z�3�9>�s�핆���M��������K=����'���m�L=�N���O��n��i���?�u��	�*�鄰��.oZw78�x�W�F�O����9�0�g|�T6��Ah�F�fO�S����8��ҿ��V@�%j�_��-~F:دK��|xa���UL�!o	9��y���/�9F��pX�7m��;����gٮ�F�G3C��H��u1���Y��&z�����1�7��� �F�{�Ԝ�K/2�q�{�dH��z*��*:j6&fTc�]���}��5���2�D4i!d�Z����9��{=Ik5��͊dLH{�8�2�>U��S��L��K�"�o��~�J��FD7뱺�`�i}}��lv
@6�,��֙u꺫[D_�b%2��^wX��ĭ��g���0�T$�;�c�I�ã%�/ +��|�5����Ǵ��#�Jh[`	�^�Ks�/�]O˷����Uk��S҉�]O�~��C'��t�p�V1��fFȋ@�r.z����5���٦�Zm3j*F�W��J���0�T1LE��ʝZ��[��LP���w����>�ߞ!ee�6G�G�H�����>h����E�J�I@�ߏ����T��r.yvU� �Yn�h�����N�.T�w�O�h'�躽C�;Zd������$a�I7�� ��9�փ�h�M�w����kv�����_��F�ARm��}��k�~ٹ�2/TD�� �)���B,���9T�1:��H�>����|S�`n��ɰp��R�������إ=�v��[��a �c3wpf�	db?�~P>q��F�*��/�%k3!���C��ڳ���=���Q��10��}
lx�V�� G³��q�[�T���3ReD�[D]�9����G>їw�c���*~ ��7
��O����������:��ⳣ�-�X�^&�PX=�����v)��$
Z��Ր9�}�b�3Yֆ.q�A&�{7B	8 :C�p�*Tnlt>�J5�K~�d�G�7�� � �ǀ#��9�%��ՄN�o�:j	�#�ci"�`�P����>��m\�n��X����a(��7�%<[,�bѩ�]���/˭��:�.��G�ꐤs�`I��٢�$���I�x �;��ᚶ�;x���+�n�fv�.s�#Yb=�q�ߞ�=�	�f0����[o��u$>-�d���o���_����QD{�� ���S.?Y�˸�k
��Ǿ�C�K��S0�j Ȉُ�mx�5��nv�B*��u�/ ���0U�Ue ��c&�:�]��7���' 3m�����Q�T*&�_��U��Ba0{'!PS�b �z5$���G��7_�b&TS�qP�љl�/�e���2}D�D{4�v*�@Ԫ0�
a�
��֒����kPϡ�x�<s�O�U��{ m�cƫ
 ��%8�N�z����x.��tLA�����X��H��9̒o�����)���F��ϓⶮ�k��ġn;Ѿ��:�iy��+��������;1��V\��'Q	��iGyb��ݩ�7�(�� p������9M�(I�<�sC�Wʮ�D)9�4Ѻ��)�n���+�5�dj� ���3_y��1qR&��́|�y�~�y[�R���j�mD��cn�텁�	��#���僇���3����jX��n.�������qO���$zh��$Cʿ����U��O�����k��g�Z�Ö
7TL&qG͹E����.��_*N�ZA�<+7�r�G��(�Lp�������EhI��$�,���u�٭��q�M[��݅�e��Z*+om/��4��g������8۾sG�"=�m�����1�ˊ�v�Zk p �:W���l�G��K#��WI��a��mi]��
]'ZS���Xh�ɨ2چ���CBj���"Ed|Yc�:W�mڱ���)����fXqr���	l�V����ƞ��v�TF	;�ì"ɹm��6����Vk$d~�Ѱ�x;bx�kM&w���RlsM�H����Ɣw�DU�m�hZfuvhY&��B`i�܁�Aq�Te�dtZ��g�����w���"��ˡa�Emz�퇸�!(��Y�y|�]v���RP�&v/��.�j������uP
�v��bT׎]X?�f���A�݊r�(o�:~[4��%���-Mn1X��A��;}�!K�Ո�{3�A.(�
�	]K�/�J����	�a	�R"Bڕ��%���Z�H�����3afJ��aM{��T�/�VC�yPVt/w|a�n;��Q�e�[R�KP}F`Q�F`���D0F��H$�[��+}6��b{�|��WQ:$�%�1�Au|.�'ͧ$b�k1�yp���v�s�*�i
���\�B`J���H���x��M�Y��,��d�@�Yn!Aw�am�َ���I�|��l���^�-��}O~C�R����
�P��9��� ��jHK�����zAŻ�i���2�3G{��@{
9��t�a��`�g��C�;u�U7�G�ꃅ�{�80���PC�¾X��Շ�s�<p���g���\�ˈ��ô�˕(aۿ��W/Qq�U����z-�e8�M=��$k\]}����y'�/�2���W	U�,��c{k�dD����oE�j@AEF�3R��NA_#P��5��n&���AG����]��7%�-���zs	4q?�}N	��T��B�Z����2��g�ٽ�@�kJXc6�k��ŕ ~���h՗�`5]V����\�%���	 hG"�|4όߕ�ru��+_ʃ��91��w��� �j�����4*˱X�9����ҐXN�X&a����ª^��^��p�c���E�"�8����P��l @tȁ�X��;�p+��:���O��rp
׿�����^+�B���|�<�n3}?��o@r�
� �P�ȴ�|l2j)z�ˠ�D��u��TQZc�����[��ꈏ]���u��<���7t=�=�Ls��O�GN�:U��|!v�W>�8*��l_�X6�n�Q��Ӹ��$wӌ�aD+���&X�<����A���\]6�f��p��1{��4A_�E�b�x+Z�/岼%�ZLSp��_�۫͟B�/ND�Ԭ�/��Z$���.�}���v��_Bǩ+k|��F�0�Q6Xc�	��q9�Qp�]�h0�3�-'���l*�`���L)���9�-XҐ�ޢo�:#�Q�}5Y�jp�1�n��~Q��K�-��v�������ni�L�C�/�n|(���'��ğQP$�G������f��&4+���l	���U~���0Ʈ:T��]碭��F��P��)�r�O%�ު����R���v6�pV���j8��'���� 6�|��^u�{ ��UB �'�m��ŭ����/�-���pMP��% b��RH ��u"UB'��y Ť��i�� O��T�C�T㷑'�>��p��r�z@�o�
����P��o���]`�D��WaCh�9*�P����"J�>��ΖK.�[�T�U��ͅ/:*���3 ����pՋ� �{�]ku6�����r�B��L�,�g�T�2��7��tY� �95Q�C2�������n�3�Ѡ��+�8�
���D�����;�¥�K���Ƈ�@z�i�mg=q��T(H�������0>L+ay�ƾ��RV�Fc�݇���>H�jiD^X�;�	#���ͭ[9O��kj��{��������0�4�w�Q�m@}1(�tz�����ێD��{��O�ꏿK��10q�z7p[���L3��Jv �XO/��^an��.<W��]FU�?�Vm�c���/{@>��]��5��;���T�/p�|'����4��q	�j�+A�F1�ݙy�?�|r��罳C�1k�2]���L짲\]:�3�Sj j���G��</|�6�b6*fF�Ё�ξ������Nn�/&����������MIk:������0nkm���m�Iv�����o��ei�F��of>��N�?�3@���}P�q��-� �	�x��(%a��'��@m���G9�NfA��+-&�Lsj�.���C ��$Ð���a�\�|�l"{�)�ǥm�G
V��MpY�r�ܮ,S),�Y� ��J�����,׶$m�I��]��V�		A������������y'_�ʐb	�Z_2q*@���a�ۆ(��4r?�ļ�N�	�����[y�5m_�Sc�*�.��CT� �gUOd�����[�g���Q�Ǔ��}���H�z���2�@	�,�]Żq����ƃ�#�܉;�K�v�_2%� �Jd�c�?dS�!���O:#�!LE�Do�3�L��ʱ�����J2.]�o�Q��8)u2���a��D);��X0�o��8JgXѤ��۳.&u��E�t�.o�É�!/,�b���ξ�npAJ,j�0A"*P�r��L�xNk<x}������a>�˖"*j���֟��q�0����8>�X�i�*˖Bojy�E�ȭ]f�w2�Zr.��ߪ�҄�PL`�i�d�s�؎��;��)��)��Ϡ��k����,Dóu#��D�}�����g�V�n��(Ɓ�{��bj��W9#K0��Z�ڕ�}6Vya��5]�	��Ὸe���9�ǔE�܅KF�t#�t���	���vu�T;,���h���9�nqQ˚Iz�
���_�g�J
FT��|j�h?�!3^.¹P���!���h����U�e�P�%�Lo�d�Z1������NP3�T���������
����:ڲڷ	[�p��pfR��8�1 �Ċ�U���sй�}�WI���ŉ��x>����]�B�L�z]~��M|�Ҭ�{����9�J)��]��X�'��a����Y�����>	�-�/%t@�e�v�,��7q�$�}�7�è��H�$,�鍇����T��1F�ڌ�(�F�<>�;�<ah�
_��bOA��¦8H!?���� �xx!�*��ۆ�XsJ����O��a�Cq��� ����}����[���$g�+�u�	f�&��v�2{�*�!�;H������,@ݻ3�2F��ۋ8�h�c���a煮��	ޒ\�k�Gz>�M���@%Kd=�	��
���(�/N���V�����Ќ���Ʌ��jt���^98:x�Y>8���(��5�5~؂*�<i��(�Y���/C�������HEq��BL�a���&$�j��b>��l��q��<�4܉��0nl�FBd�؎����s1b'�R �����#�ݷ�����S3cG����k�F%=i�{�_x��S/(�o�z�vZn��Ļ 9h�$M��3	�>c���$�B8p��T�'��!��|ZJ��+�� �Q��D���*_�/�esP�1�`�*���%nhݺ��k�H2�Fm�G���t�6�R�|��_�^�}z��a^IQ�<�Xb���B��b��ђ��AO	�K�� S
�'ih���,@i&�^�ۂo�bmv�eTJ���X$��X��Қ��G�rh��7E��2�d�������(�i(R)/���1e�E^ؘ��(�bd�^t�[O�ٔ�P��X3�.��~v|2��67$3l>�"�1t�y���׫�^��)�T/wn�&�)Uy�&!=�W�S�bl��P�1�NQ��yx���r\��K��vOw[��>B�".'�)"�^�;� @�+�.��G�i�����4F�j�:�2|�>���߀wJ^'�Q[�tA���}>�Y��/V&ul���;2X���jRa<�fR��D�Z-ˆ,�?�3�Թ�o�o�Ч�?if��qr˿{���=62�~�U�p0���0�L�n��q�T���!DLB�_]m_�]>I�#�W�fĳ��'^a��$}k�E2��ܱ�ӻQ�"J�ÏD<;��4�Ν�	sz�+ I��.�R�<[[BL�<?<F}By��v�IX%w���ɀ��%N�0���<�	��7�a]���J�$�pd-HG�� '�����J*#�����&��O�%��K�� 1�,j����:h��9T�څP����Ш����1��z�~�Czb�g�t�4��%b_��W,ZhC��m�2͋�i�C���G1��/�,��D�6�l�U���R����C�c#�y�Fv�bB
��Y� `�6�c��2� Y:<Ψ�`��� ���HԘQ6����k���4�]��B;ұ���NC�;޲v�w^oѝ��Z�o}|u��C|��6.5+!>@�5���7�$�f������.���6כp�P��<�ђ�'�N�ܺv9���À��|9K�L!��ڽ�ջr'�Q�g �B_�@�o�HE����jo�-���z�R�ۓ��!�Ue�;FT��jb��'�Z��ɯۆ���hL�v�/"��ec��eu�u�q�^�:�A!�s��9�fL-S��4\�X�hm��ۦ�$Z�,���nB����~R5u�j�1:O�.�Lj3'�}ϐuob�zA�$VPp>�|g�?�jm|?֚QaM'��~P�s%��\�j�uAW��^�>��y4W���<��L�^� �`3�#oy�%r��]s �0V��O���>	<Ⲭ�\�I���/����JQJ�/��_��:��R84�+0���N��Ŀ��i��1Щv��	���pDO�8��uoһ�˅�H��e`D_�M>�4ڈ���WNV��Zj"�+s<���4�o~��b�!��4ܢ�t��sof��e��o9�5�֒[�w��%8T�A�&���X�;�\�P#
�qNf����ѹ2���\��/w�qW��w�	�w�C$Ѩ��a�]��
:�9Y����楩r�g�d���5A�L���R��DPk-����\����^/9�P-����U�+�8�20�j�Y"�Cpɖ��Jq)
��^fWo�&�bn���"�Zf���@h�6ǻp_7G�� �w2�%�K6L<�1�f55���,�=��`1��N�C6c��աϳa�/<'w�g�Z�����l�z*�������V�&�+c�>L�Z��b�nYka�H��$<. 2��m�k��43�b�a�2i��UyR~�9s"(�E2����*�F�{�?�X��8?�����8,�+��	w�	��i&�aܣ6s^�oV@�,0��y��l�lpf�s�
u�!q�r�^����M���(B*�Ӆ? �,�`0Y���?e}+e��/��*�[��.A���Nv�Efc@{���u>f
x���c"H{��/����������m�ʶl�2���nq��)�* vAÄ�IH��6���:�Ot�n�����aN�Y���?�k)~�lnHxү�Ç���0
n.���߫y^ hsb&�������M",9��m����v��&��LJ��7ASF��A()�;�";�Vㅔ�)�ߒ��P>�vm5��Q1Z�c9|���`��y8��ر&7��4���>��!���}X��K.�p
��YwX���5��Hעo�(6����/z���5�G\�Pw���bc����Ҫ���� ?��RŘ�@#Gh/f���\�xt4��>����\\K���uK o�X�� �{?z:V�p2n����<~�D���$���J~�ɂ}N��U�n�3�`{��k�ť���9ܮ��0*ُ��O�%���#N�j[=�^��5��}�ѹ�-��N읎���	�^~Z*>.����\ 5�ya@�Av��?�U˰�3�C�Oxy�E�k�zvG��M�⊨p'8��Qa��1~ӂ�Pal�˪�Z������e$Gv��~-�)�G������}��詏
P|��f���+�
�t��$�͍��A �$0^�������'�2J�Kd���O�3�a�QN�� ��V�o�c�h�x���P��~K��L�����ݥ�yV��?H'��b8���B���:�=���ߓ1��ϭK�ʝc!�'x	-���7_�[����0���D7r���!s>��)¦���ʭ�>?�L��c(y;�`�f`�G*�Bk�Ǉ-���FR�L1������B��Or|_7��#���>�F-�X_u?	���i���VtL@�g;�d;�Ӽ��	#�/��S�ąr�$my�B8�miV ��r�����)j�׺]F�AFCa�x��B�2ô\��`+r�������k�نl6�o魞|�O]98T%P�$��ǆ`��	h�f�E�E�:'�����Qķ�<R�thgN1|!��:����krvk��<E2!ޠ/�1���2�� 6:hs���O�`$����^� e/{�(���� �n�uR�oH[�^��%M�mM��)=ճ�ف���8��Z����	}���T����>|�9�����v'4�`P�ɛ��z�Qr�X&z󠎶�;@��=��#{1���"E����y�,�@�E|#c`��B4L� F���J�L ��}�����Gm��5r:��C�Z�/X@���#�R�@5�;�������	�1X��BҼ��o�TNn�<?��-��r���Q�^�6���SQ�a�,B�ˮ�R ��1?��ՠ���PVӉ��+��V�r�k�"f����v>���p�~"��.��?��T,9���2��Ap�eTg��@��d|�NI��=0�jՐ|�a��pfZ�@7��T�(y����#������=� �Z��I����eo��7��X�ǩ��(ۼH��<�R�B����+#H�Ά����^˸���������tԈB���,�㒝!ٿ!Z��M�m�Fa1�L�Պ�18��C�7�3���J�oGp���C;��Kcw�� M�������OvbG=���Ɏ[��?6�ćI�;@)"�&�Xwz�4��,���j)a��}�U/���JQ��"�ؓ���0J<�Ma�߁N�r2���U=��Rc�Z��Ǻ���� �x�����$����.���Es�viT>�|�B4_SL�lꎆ�@\�г���=-�#EWxI{��}�]Q1:UPj�A9ŝ�������TօI 5����ӎ�ɀ{��[�Y�k�_�����i�8�D�]pV����O�濓5���t�.	���_��;���Z2i����K�u3Y�HhfL�砛�?F��j#wI��-��r�h���N�в�v=�H�����ZoF��ڶ%K#��p46���B%7v�|u>���ӠhR�gJ4W�9΍{{>©Yğ�3��k�وH����D�!t�~E�:�o{�E����0�1�����v��M:X'�D���|�i�sXƀ6�o��D��h�5u���JE7<�p�k��4}�ޛ�Ց���f�5n��"�u�r��R��6���i)�~�W�Ӏ��& =ܦY.�����/P�x��5����Td���;��!h�s^��>�ړ�B� +�I��Г>�P�A�6��W�/W�*\+��8��j��!�X�P�ge
r����`Q�:�H5w�[Cĭ�=�qQw��N,��ؼׇ6�4�]%���DduE�iB��60s@����\'��B��	$|���k�K��.�;�m�Z:E����:����F|��x�3�8lf�lo���Y�.Э�´�W�5ado|��֔��ҟd��*�+�|���Ⱦ+U875 ɮ"�~�9%��t�˿0RY~,�z)�f �a	�c*�
�hٮ�~˾?a(P�����d�i��k7q�'�� |=�����`��Z^Fv+g%/�1�੘9p���M1[g&��\��y�QT��U���z����_y�lfK�s�J����8�)s�!)�A�2}��2���"�: ���T}��m�x��o�������k�x�b �=D)����:���ih5`��7�"u���H P��+ﴬ/?�'�|HǴ<xv�	o�{̃�%FG��u���v��3������j�&�{��+Bv�\e0@����cHᾕ��TCkɍ\e�sV��6)��bʮn�rç�BO��/l��b�+�>3q�3r�I��˭r�#dƍ��.X��������P�J�� z+[�
k5M�N���"`�ZeK�\!�D�]���-"s�7@����u��+���5J\��I�ݔ2��C`s�ڬ1�㍐���fDt3�L���ZIl]�j�Pl���[��$���_����+؄��tTt�-�d�ڃSG�eoQ-��TP�N���8HN=���Ă�ç
�F<+����2[=C���t��:�܁q�o�����h5'����$𨧮{���;#h�`���/�m^��(�_Ĩ�-���ߚ*$Q�a��r�#�*q��#��N�����t�E������t�K�,x�t���dB�N�vTu@:M�9��q9�l4�q*�EAn��T��pȄ\kF�^� ���ְ����! =k�������-�.��ru����s���=�7�a>�&5���"�K 5r�Htv{�m��*��v7 �R
��Ѝ��q����dA���^�F���С�4�'P�DH�0D���^�h���Ky�?B��)-������H��xUX��P�y�鋒ZW@��M���j�
��k>@��_�
l������&��G�y��Q���E��q鋖D�؁�^���*�ҵ��c�[���t�۰��'2Y�s���>�Mq�91�����d�b�T��0�X���9�>�4�������Pm�LM�謫�����i7��;� Tշ�sh��u ]�(Ho���Ϳ兽�c���RW��~���S��� ��)Τ5�;J��U��F(;-{��L����r�z91.�M��`������j	�~�D1���C1�i7!��(�\h��l��J�H�-��&��:DD-l�v��S�EM��l��U$��Jr;�Rv�Uk�-�,ø-Cr�>N{��?vU��G�M�S[˶�<��EGop?^��x{"�R�/2��ۻ���ｨ�|�j��IahX�����#��E��M�P��������J��|���lr� `�� ��m�6�X��$�
�,�0�.����B-������t~���M���HF��!g�0첂�9�.F�����p�f3���J��q�)V0ṳ��U�k��С?�'1��3��ڲPz�zBlH�K\��5�J[]T��?��r`�,��l��Z�����REZAU�>G�}�p��QU�\��u�|+(N\��Ԟ�yk��!�㏥y,��Z�^�H"��{�^e�� ������)R�04�����Y��P��`a�!,�T�R�fBYЌ�,��p��]���v�T�>��P1�1��\Jކ_��ϔj��V��@$�u'�O üf��_v5S)k���3�Q�C_�J398����>o��1^�30	�b�*k���?1q������A�P�淉PUT��e��v>X�_��E������)�����&`�A��C�Q"#Z�>Ky����{�ѷ��܂�L�H���.��0VX�3H�Y�@���ou2,�qqO2�^�$n����/\�=��t#��K2�s����և�������.���������ς�"W�vhW}�C��P�f�y���v94xL�m]�c����v?2e�F`��
%'��6�������R�P
>!A���7��f��C�@q��k{���f����b��f�K)B+�(�M�	��ܘ��;H�p�l�L�|[��E�<�5��Vf�I!���ٱ]E��̦�T�U���"R�1����9����� \�'G��Ծ��1�95�?ej���xR;����;����D6��.Ÿ�c�i�I���T#��t@�X�uyTV.SB���N/�:�[.�z����	�÷k"�����C�g=�?k�c߇�Z���ҒO�~`��~�_���#��6�("՞Tn�O��L𷕫�l8��$���ť���C�D�Ò��άFN�;3YC<��Q�k��w�_��2T�n%��C�^
��m.��T�/4�Ŋ{
f)G�T�kZ��^Z��AF^�W/�"e؜5�b@ �Y�=2�AtãÝ��*�Sz���0=�y�e�nTǓYP�q�"��)�v���z]��#�=A]��䐝��<�QJ*���A#�$`P���"1E���|}^���YA�Rz8��)��k��\�~�儿"NB9{��`2rL}H	���A�2wa�<�����>=�/vd���	$�����4I�O�2�+�	�X��T�tt��lQ*�0լ8�6�0�o�%m����&�ܓ| N���/Y�|����;Ć٤����ؽ�haJI�6�e����=��қ��T�	K NwP��"�����������E��Y�Ǜ�9�kB��O���y2���9��O ��T9�R�@��5e�|xLq��4U=�KJ�/'C?`�Ei>��h��(Udb[�=�N) ���j��Jt6�~�G��T�r���=Vp�����ʄ��0��y�'}���30�����@�A�mG\�]�0vFZ��#C�����������N��e�빺�qֵa�@R�br�&̈BS+���ퟌ��+��н_ž;�^W�<0�dc�ԡH���60b���.���X$~�,�P�%�ŘO3��m�2��r��2��e����!�M�V��'�
H��Cp�$������pBz�����@(c��s��z��a�^�\{$�Rd����w7J�9쿇�.A#���������!V_X��.m�'� ^����'ml|���@�O�r[>��|C�/�φ���c�|��A������Y&e��8]��{Fţ�Υ�_�>GHo<�5lfd��L/�uT��p�O1�]�`��T���z1��X��ݕ����Cp&��'ʺ�F��)��^s����&L+��^XwT9k�S0Y�WAGn���*u nW��7R���.ߋ�(+)g�(�
	�L��G���@5?a���Y'��ɸ��f3�rE� ��Y�@kN޺�x�U���|�޿9�?�H�{�3���[r�A*�`�P����\�ݰ�o3R�H$+�r�<e�"n�8����K�'+��=N�:�9�u&����hT���U�J����xaN�%?�(Z�;\�(/�=��ݐ���j���x�9��$9+<���Yi�G8�X�$pR�����\\�b43�B"L����')㋟�,�-r��;�4\A^l~�1
b������P4�A��Jsx�SCg4]Hu9�q4�I�-a�cʀHH����j�j���j}�]/4����ڿ�#�h�fJh�/��PJ�9�sG��M�e=�<�嚼rw����\F�!>ZdѢYY��~}f=���<�u����Ѥ��5C	j�����~�J���n�[G���ڠX(F!*�C�E-�[+��u_�tס��YeU�ޚ�pž�4��A~n]����Ze��̕'Ģ���z�Kl�eU,����i�쨾��R�,�Kl(�ms]�U��9 ��Qُ�j�.�1�+i$�Ai�sm���~I4�ʦ�}�eD�>�ك weq��$ڹ��zV��T�U�����R�>B�3��˲�$��#�4�\H�.�&��:�����׬��8F����8R�'D�>���g����q�M=�sn%b4�&�,�]Eϵ茵M~mL;  �0?�y�ky���8����(+o�7��I�ǽ�����e�UC�T��_��]�u0T���@��;Wk'����eJ�c~ݞ�e�hT��]&Z�o@BsEg�'4V?���X8��q�=,3��*����2�BϬ�A�a�����ӿ�ѽ��!㼼�U�~���DwFq0���f�iH�O>��<u?��\��q8w�[��[ ���Դ��pD�N�{b0�/�sΗ'�V���S��,��m��-�oc��g�ˇ�
��EL�����3�x���T<f&ϣ�ɫ"]���_ĩQV�t�yk��ϊ���d@��x�&��I���Ez��ඈ�(�|�W���Om<d����� Ɲ}�#cC�:ɜ.s"�6M@ڛ8�Ik�{�󱧓30	�+������M�M���������hi��8����b�y͓%P�D?���<.�i��(�V�%��j�v[�b�lZ�p��W� Xofbz(3���\�P��'yJE	 ���2�����.TC��|�%�jpe��۞���`)d�UlC<�
��������VBEϿ��CAf R�l;����+�ÁH8ċ��1v{N7�Ndv��mw�r��q�h�����7Ug���>��
ykT�_�WC��f���Mh�����f�ͱ�:��N� B�j����헎��������u������	�X{Y���aD�RG� r��2z�����M��~�2�Qm���2���@N����c;��%^���տ���K�
�V~�~�n0����|�0�u~|�_�>EZ����92o�U�;�2�a�犯e-Ӥ��� QG9W5��7������d�eHJ�:Я],Z�I\fQ���]��_"B -ٓP�2r*�8ǆ?�qƍ@�a�e�|_��1���M�ð;!��T=��ĆgU��}��i!}�i��_���Z��0��4JT����0���0"�/HVz�䁦ɼ�C.a;�ټ��=�$�qط����.T��L��T�In�~��m�߷e����E��8���p��Ј/�`�c;�h}�0y�(	�י���AK(-�m�Oa8����C��7D�C�X}J�A֠�b��ue����Z̀�Ȓi�M�ƈ.Q�ѥ����Y2�n7c�ӳ�����W������Y#�Q�3��	�d�\Fp�L����tMJ]��c�T�������E�(iuD5ѕ������/����Q�7��͹���[W ̈�~Q��̍�N��LLrntڐ�1�$��b��j�p�")��9�Υ�Ɉ���3�4����½�Yg��X6f�q�)�Z������"��A#g�i��{/(�X�h��7,]�S���������|�<�cb`Owz���,+_%�q�9H^���x���w'�ʖ ���M`�5��3����S���8�!�a��\;���)�B���(��:^�SI�����*X]]��?��u6�<� ��T�����7��)�rYao�DH��/Ψs�!���u��:�ȈG�ވ.�?A���v�FG�������/寧>V�e����V_��x�z�[��?�{9QU>D�޽D��1[2����P��N����j_�6	��>�e��]�pɶ�':�U��9���J:���4ok�������Q��5�zO<��7���m�P��rWy�T̷_�+��:b���?(v�7��{\����. !�.�3z;Ԃ���bB�ݯ*����H%�O�d�	��k��vA������s�����F[U�8ݕyu3����,o3��A��޾r�K����[��:��xg`}O(���`-^d��aD���R���>�C^%�(�!�Ʃ����Z8�XA�b<�����pa�IL�����*�t�\�*󱷎�քw���\8���XKf�o������J�7�.�Ph����G��(���_�!+Ԅ�
4!�45�ퟄ3@�5w�"��!A�p�m����l���?�Yc-ֲ:)w!����ym��s�?R�y��H�c�)�Ά��թ~��і�isV`~8�˖l� >������_v,K��x����]���2>;n������4tG�w1�e��{����C��1͇hξ.`��C�h�K���xΣ�[KI��C��q��*a�s0�֤]���O$w���-��.�9����_�J�Zj
��]�LM;��q���d�լ�r
����������=A�L�{(���!����f��f31�0�Ϯ���J
�?���hדRʏ+Ћ�>�r�H��L�ڋ�ԄΩ��� >�kVNΥ��_\�S�t�HOה�<K�z#�n�Ԕ�= �}?�ɬK����X��8*	��5gk)@�l��@]���%~��E3��n�7���v9:�􏎁o�{`���Ć���c�����e!+��?ך/����P���ŧ�rĒ�K��O������c�q��k�_��8J5N�$nTL���$�ۤ6������v
L����h��U]n&d��p#«.�tGNU�����"�dظ{D�W�5��^��ZHq�����B�\$m��d�-`ggԼɽ-��Ra���h��{c�J�Z�	�_]a_i����-ʙ{H�$��'�-��ɸ+w�s��B9���M��W�.1�j$z3�����Rx�'��v�=L�?	~V�by������w�"}flH���X�WC;�b�go[���Q��A�x��҆�H/��z^>lD9���ݹ��8.[^��ϙ8�_� �t�@�p�yP�"]��G4ʥr�#,.SlWF�k`�]�aV�
_�O"�e��0���s=�����U̻��SZ��C��{se�KXt��P��� �Q�=f�BC߈�y�󷫴�Ws�z�Z[3���ŏ~V�EQ��ǉ��0�����CY�\8�-YU��jx�Ⱦ_�h�7��F���q�%��L�E�$�'U�%y"�O�����$���x��)yGH/Y�s��N�G:AJ".��oFꁯ�2M�Pe)��(*3�o���cT�w]�@�鍂�&�oj���`NqfΝ߃�%�%�����VI��I�VeP1T
�+W<��[eȏ��KrD�֗E�	s:����2S�VL@��l<�P`� )6�S{i�u�O��,�0��̡j���"��9� �$e$9����1����"��3΃�)˘���E��\? |�"k��,�:mu���ȕ�:d��J��A��ș���M���`�ia�����N#��.�xE�l#)�;���ͫ\��q�'�2ZFC�u��K0���+���XԼ\ޮ9�Dc�W���,����p>�9���<SXh�2��_�"���}L�S�X��ԃ.���{x��ʉ�IN�Q=RH,�Vi�C.���L���sG�h����։�`�����H̸��m-REM��պ|'.�K�b`�(�+`����~y��4�5,�i��?8{x��;�Z??��0��s�ϪxZV��^{�mݥ��yڰ�6��bw5�䍲�������ռ�TR��w��W,S������x��1���A2����4z�Eİ�rYF��W�+W��;U��}+<��Ij/Ж��� FO���&�V{�����������j�S��4@�B��8�����=C8[�3�� �{����|Ԟϩ�=��'��I�Yr ;���:��#Ɏ��G��E%�x�`��� .	�� '�F�=
D���`�A��y�������c��}1�)��8=�US������>�7���ǭW�?��@X���b�k��܍�Ǩ�o�4�����߼9#��H������  ޝ�,��lfm�Y>Q�i���`k7�$$��d/��/�$�ot�Į��L���������#����:�ޙ�S��oO��`lS���Ԡ-@|��pۈ!�t�!&m������X��6Es�#���ڙ����o2�(�LnŅB+��)X�vU�#�b�H��<��З�?q�O:cb+�9����7�_{(�f�ڮ��b�c�p�����
WQ�IB���@��j��[y�"�+��$^�y{��B*�6&�ź	�ǲs�Y�(��=�9= A�P�ޓaM4$Y���X�KIa���d����Rn����>q�i�h�Djn�ۿ*+��,��jn��Ӓ�&�p����M�j��_���eQ�!��B_�+��I���s	�q�~BQ��O�2<�n���g��#��LP�C���A��D���)��t��3��6��nMO�B�Emc�����(��|�i�!ǃ�t)`�4%��4�C��[���䪅�
[�^2#ud�K@:{���ee�o�D,E����)\k������ygf�6AyG��Cr�k��[J�*o���MS��\cqQ�2���;"\j�h���"�5�N;�vF1�������<���e uZ�9�N��[1��Q[�[�|4c%)P��-aE��,Sp��Ժ̑�j۰�F<�]ٻ�V*z�ׂ09�^�J��w=M䈲
�����l=���}^wU�K�Ũh]&�?�)+�=2J6hX�	�����񳑡ۍ����l���x�7:,x��h����(�J�5�ǢlV�Qa�ȰL�W<����dp��
��g����]�������;��`]��>�<��($Y��%4#)��D������Ȼ���#�࿁��X�K��f8<R-�R�l+}N�m�ܥ���A&3?�U�azO��Y&lR�tܞ��uqNE�������&��G&n�,�)VBퟹ8�$A�	��r\5� {��<7cz`���;Z��Kb��{���v�s�d�J*�")��5�Y�<�����,d��zɜ6H��9!�^��ebԳ��OzEاTC!��П�!S��ӳ�����kt����MZ1i��r������$���S4��y�x-U�ո��z�`�|�B�F#rQ8��q��qr��K8GL-VϰR��������d �X[�+���wM��n�>��W�����$Ȃ�U��/�ZpX�Ѽ䢤�
Sÿ#s!(��RX� FPv,��@ "q9>��:XY�.��"�IS�e���⭁�5_�U�9����(;��`ȶ�b�u�}��01cT}T����W���44�'����D�)6�ci�%ѿ��M�%S�@"߻X�^N�E}XS�(4�/�Ɛ�%V�ey$���uVx	 �Pk�Q���)��y��V�W�)Tr"��'�@��ߒ�vX+����v
^-�Лĉw�
R�(��
�E$��g���� m��`�T�E"K���`�Gq�J��w,���>b*ڽ;Ȝ��9^s��-���g^nR�T���Zn���� ������{��Eg"BJA�]���f'��)<��v��͞���'�CŦ���������dbx�dױ��Mr=n�3e��=E8L�1R�#�4���
>g�l���M9.+J��nZN��nm�T�D�n��;���N��3��������BkrUMj�g���/�<݊�Q�^ї�f��t��:(7`�Z
U��Ŭ�ڬ��>���� X|�>�u=@��dhD��������u�M�s�`+��qM�Z�:��D�k}��֐Iόjfxd�U��uC�dQ9Yϡe[-��cۢ�D/�G���Т���>��uҗ�s����#Й��NI��/Hv�	<
*JOcN�:�ݸ�����B��������䰅���m^��c�e�j�i�]���!�gY�F���I�e��I�-3c�GSm�2���O{fkTOq@3U�q*���f{ �UT������� "�{����߸�%�h��t?"e[�@0�,���GO�o���M����>�x���s-�^���u/~=�v)���\{��tP�,��xJ���p����}���8�u7ƻ"��8ya/�Z�\r3���ǡx�>�x�������*X��xc_�Ϗ-�4�v������?5J�ˏbx��fj����`���pol��4�"BG^,��sJ�[��p��z<�|Y�S+���2p%����f�?���<�p�Q 峻��진����t�:Ш"&q�Wĺ
Cg2����)�S�So�#���}���5I�y�:>̾��6��}Ջ���NR6��%�>ؠj��=�K5���(y�sctҞz:%�:�$���NP���I<���Cܷ�0�d��Ъ1KjT6�9a�(�&�Ӵd���6 ��L�`���-Ro1�yi��=���#gP��l[c�֕	���3�#~����2!ږ�oe0N�h����e�I�5`��[x-vnX�a�����=��bj��� ���j���¿2v��y=�b96������#n�f��d�ߎT(�^�R��"Yr\�1�2��ڄ��_��_���{��SV��ߡoN�0ԙ��klCYdI��?|�v4}�w�@_�����3�(<%ds|ibEt�����|I�J�S.�	��eZ��\����s�/����v��$��BQj�����V��[[�w��y���?��M?�xx���ҩ����5av�Q���R�;M�}.��]��K���pP��-�p\\�+�ݬWY:�$?��K�As�d�1DóO�^�h�^�1-�<���¦�����¶��:�>��w�l���s#���P��6l�D���d�!Y���o��%�LVްvC�c�������@?���=wQ���Ť�Y�j��'3!>ta��Y�_�9X%K�ҕu�X�����5OQ��O-;���ٻ�:)j�J=s+g�U9@���S3=M��Un�9?�.Vr�ۯX9&�������v�|?2]Km�_�|��z�Ԋ* ��(4z�9�)x�1�jK���^�ú��X���������;oH
�鏾�-����T���XS<����ɀ>�5(��NVU�{d����=S�NQaq�7V�]��y�W��>�aؤ��E��)��:�r{D�ޞ���&��^m�e9�^5;���xpD���qte����XSv�/9{�"�nG(
��He��h�'`qǩ����k.�N�����w4u�养Ey#���h^�]iёn�U�v�;B���x�*Ϫ���ZNVu�u���#lj�O���Iܠ���RM������v��$���븤�r� m�+�.���k�MH�#-�%Bѻk50��?���uu�zT�"�J������]��U$LD�]��ƕylz�aG�M����e�O�j#I嬌Dq�f�*�Ԩ\ƀ�o�)E�3�h;J��@l���8����n�R &����������r��ZԧX�]�<'Q�-��j1#~�L���>�"�<�v�{��m9�I�f��a���|�n��hc���h�Nޝ6��#�5��TJcl��g�c�B�:�E�v���1 Ti�JP�ʧU��[~��O�P����_�x1w�E�K"�iII��f5���T}���Da{��bd�wDQd)�X��쫆��c�uFX��l��-6IĨ���o�F%��`� �\�aP!41դ�d�Ę2��� ���Hd7�RA.�D��t��I `ǚ;��}���V�9;�O��y"�k�Q����w�pG��9��T�A�R�7'�2�x����sE9�s�����7M�?�,J���Ln5�MW���kl|y�o�ê'���'QZ㫷���k�i�3G�J��m�4FA��J�� `�a�쐻k'/��^�Ǖ��׾�H��i=�[!9wE۴�q����V��v��߂���>&��Kk���!��o%�$���R��M��3�LE���E���~1�y�+�sw�`�ZÎ��>����	����nE�܆md���Dms��~x{�}o`��E���������Y�[k�梍�~W�ѫ�}��2�4�+	c�������h赡ť���9����_��-u�ʬ���̔}t=�Bm�Q����,�
��V��-#�Q���Q��zw�lO=� ���zfc=���(��޿�����_q�pї۞l�p3��+�5�v�ӹ���ж�Q���ϼ&�W'i��gj��Pw���0�߅x��ݚ��<j5���2*����t��'y2lz^̭oᯌ�HwQc�{1(�"�$xCD���.߇�$��4�#��H;�B 1���㴤��U8�~+[T������`�_�Q�d{�ʣ��V�g�W�8��Ս���ޗ���ә=+}��ED�5Hs�UIN\��f��]�TF��9c�~��<�m@!������몞S�Ӏ?�|a]xܿ9Ni�<&]B�c	6X������(�u�K���4�
a5����� 㜁�6+�`�e�X�bΠ�R��(�� ���s���8-�Ҧ��Cྉ��歯X�,������B�����W��%�W��RT�r��Q,������܏��{ʚnq�1�HljW�l��pv��4�#��P;�K���1,��&V�.{��M�_����u�yM7�6r���!>Ny\K;^D}_��k,�s��)�X��!i�5���L�d���B�1x�I�}�2z�����5�[M���a��W���*��t9����᨝����X=j^�T��`r���`"���YJ��d5|�<���^�Ǯ�Q->εCu��]g��>^���"����J셯z��3��Tp8����v-�k9�ߒ��6��׊�|)^ty��&(�����	���[�U[mS�I��BٞQ(��h6J{M���PL�YS�r'�ǝK�t�#�K<���%j·IB�������4q�n�߮���t�/~��
�J�Lz:�o��O�m*gs�B�����=r�H �*�&PD"����4�к�7[�tdo7DO�U�% ���P�?Bs��+��X���%c
o�.�z��g�~7���4��LI ��xl�6�e�m�ie ���R�C�h^y�������uσ}j��dpp��>��&9Vt��`o�<�TO-K�(6�zO��Vѷ���#�9J�h���c�U����,�mh��al*o�mn���>K�=1��X����"������*?�zzng�pϒ���,��7O�����$Cn�* m��� �kwN�48�D��㡵�����d�QX�6,�}���F�p������:Y�����ZRB�N�[:Hz74r�)��gB|A�*e�NZ�@~*wR�_������H�7�m�P���7��]"%K��~��M�.-���	
�Wp��6ڶi�t�.~WuGi�s�U}�uS�*'}��^�/�/��]�vE�*�ޜJϡ���M>�⢶/�r*��>v_i%�Ds
��.w2aYp`�_���|�kDA��ʄ���mr�������ʣ���X�����=K�f	��Zw&��}����������&[�~�������������B�3��<%��"-D���P�ta}���pE��sB�[L�d���JT�1ֲF<GA�\��)��΅�eY��eJŅP����!L��W$O��֘�,&EV�����?\��hA��AY��VQ�w%
�z0���D`��mP;`�~�­��$]��	Ǥ���N:)�E&�`��!�U��5\~�ǯ���+j��ȷ��y��B,ȰC!�M&�J$܄V�F����o����k����|M�Ӛ���g���a����t�9���p�h�U����[2xEJ�	�[++�=��M�1p�E����I����Vf����ce����]��;��m�K�~AMO5���nL�I����E�Z�e��l���ڊdGs���#���!����w��dM�iBi���7��O�%�U5���Z+��<��̟�IaP����kM�fH�!�ư���� ��1|�xM�vY������GU�'�p�!C�a�z��6V���YΫ��!���x!��i�	3��?I`��;Db���,eO�*K�Q��|2o6�f1qH"��G}�
��(�Ё���q�/��-%�?��/-�NoBwW�:��]^b���B���T��n����󧨪 �iC�w�/8�5S��U��l[s���_y2��ƥ��.قZ����{���g���\�GK��ɷM�&pg>����H��XV��>/DIA,���\DG�R��Ħ��KzUM���]PH�<d�ᛸ���E�X��Gx�L|�Yu���m�����G��P�S����w	�q���c�{���$̌=Ђ��������¸�k��q�Q�(ʽt c|�C*�kR��b}�H���%n/��T�G��������b	��DF J+¦	�h��3����0��n%�N�~�\�;��x���X j���JM��rb?�z+>s������8{t��HD���8���T
�����|��
�M#�O2�7\�b\E΋�D�ы~�a��߾�A1����6���x��Ӳ����u�ˈn���1˫eJ�B��15������`���`�����lڵM�"S�
�6K7z�����[�����A�yw4�Z����vg� 0;�	w��mcw�r��	>Dv�E�Aa�~��W�xu�2���|:ٰMtk���өۯ�S͒��^��o	{�L���օ�f��4C�]�6�J��R�2������Z���KrWaP��`ʷf��0F��p�7@EG�je%L��W�М �ƫ�tH�C'|����������AU(p�r��������}0F�&:��0���K�\�l�p�o>f(w6,dU=���9Aa�&�&dR�n�F��C��5�Uٰ�tb"�2�����Ha9kq�bK�}Qj���ÁP���Q�*�y-{�Y�)��v�踻e�<|I�!�w���PM�vV)o"��{�PN�<�U���f�E��e�͸А�~�id���%���n`Z{˿�9C����+A���^�0��!Vމ�k�}��dQ!0'�	nHqس|Ӱ��j]/h��.�Y��4����Df��������u��[f8��┛��i쳉)z_՜�M������:�I���_I}��g̒��L}�gοm`�q�Ȅ~>h����C�n��i�G����H�՞�ϳ�.��:���^���@P	F����}G���.^	׾ ����O�u���L���{���V����E��W�����`�E�A=�I,i�Yj�ԇ~B�76p]E~���<I#�*[�_�*������g��}N6��iw�_==
4��`�PM�m��]T+�2;L��9J���g	��ȧm�L�z��{�Ms���S�s�G�JHin,��1j�����b���jVNP��i5�T@	~ze���͈ ���zXN����a��[A-�˨$)��W���޻�QpV����nz���T���<Ԙ�KOU޴
\k�����$���}��y�8�g|�2��=�,��	�H�S�b��T���k��īX1�C����ED$�l�0	(vU���,�nG�|B	ih��~�Nʴ��+�ςGP������4O?�d	���Ƙ��\ϥJwOB@�H@�#ɭ�?�D�phy937<@��p�:�����Y(�*�[c'�t�$�αx�0��BU�����X��=m��0
,8 �i�F��ʟ����+�Ja_�{
?iG��ڃ4�A�}"��C���@���%�����0Ɓ0;����`D�$�0
pozu73����y��Kj�=ݓ�GD� Kzz��5�.����W"�Oi�ňnq��׸�~o��%Wb�h8�� �0p�mPO���d��k��Z'�WV��6a�}��a�H�j3z�̈́S��p��y��5+��j�(tdl�~4�3���v��3�� 	��-3�VE����ﳸ� ��<��1jצ�\�G�=J7�N5]��l7���ʗzg�Q�m������Z�|	�&�Cp��%BGj4����_#IX�󥋊Z�<�~\OD�"Ku���E�P���9]�'B7��-��7���}/�G�����q,^\
܉���)c��'W[��dVD�"�<&A�=�Itz<�!e�o���~,o�� c�76|�,&�� r��cx41�@"�W�}�-&�E��'4�4�2Q�]$���%|�7��羪:X�}l��7�e�F���1��ʸ���Z�m��C�
s���a1��_+]��aI��w5���"ޒv��ȕ�����;��.�{���Tr�;��������������3���ZVu|<8Ř�Z��2���R�w�Df��&���,�Wz��[OU���Z���xQ��L����� ̾�oy~<PH�]~�GA�U����w���e��N�i�aW|GF#�B�c�Ȳp�� txw��F4�-� �g��X�Q�K*��LL�o�~k��<OA��D�Hhw�K�'�����^�e��o��r���1����I�[��˸�sb�|>D�/p+Ϳ�u����J����^�6YEdd̓�WkР�+1��Z��oMЊc�f��[>��k���)|^C�-F��C���n�߈'�`Ϳo�!Lų������	`���Ʊ�K#BI�k@�{�:B+��p���1�}TY1�πMWf�EwދA��(��m��d����t�q�%/��\�ջ�9��J��Y��R��VC�_��e㙾t����S[`v��b.�{5�xr8Ar�K��6�#�)TS�G����7�E�Nd��t�g{�g���1�����}�,���Qy	�ś5ž�w��#��ٷn�$��񮖺��oV�`2M��O��s�kn4�F������H#[�и����R�Ȫ�����JDg^���޸6EAx��-Qf���n�����љ�'0f�`;~7�}n�������I	��g�`˪YĪ9�Ր)�:^E��U<��L(�}v/m	�Gΐ���>I�+���I�^�Vb.�� S����O���Eղ僑HN��Pc҆/�� �\��[��n.O�a�h�p,3!� Hk25~�9%�M�����DKN��YB۴SYq5�ZA;��.����х��E �������ݖ3#g"�z��~g��g�#{hdc��#L�BtaQ�W�b�o.�Dk���sy9ˇԏ���#��|iǬ:hm�g��8B�N0�ьYV  �+U5��k�w=�i<h����<�z �zs����I�kݑWƳй2b#�܊x=|�4�G�Y�.+����,	��}�*|�!'����j���\�xg]�^���Z)�{�������hO਋:&c��
�d��}��\���ЂO��z���3]v2��p�ˆ��q����6q��ޏ@ ��k�[��'��S��h̹H|;@%L����M#����Q2;����^��6�rk��Y;E���٣��#�Η�#��e�;n'L�6��&��j�wb�I�c*�̭.��P�x�R U9ĕ��������bjݨ?��4[{�y#���}��[l��x$CJ8G{J��+9@?�V���*D]X�3����$v�@�ђiT)O꼇��){����±�1��Y�G�"2��Z��B:�I�J0�RV�bn��х�gbK�P��n����I�J�SK �1���):�H����zN�Yw2�K�C��o���o��ȿk�����/M�O��OI:nʽ�˚
��+�٭����ұ���C��d����g&Zmֈ�����2j��3=m��r���qGM��uOf٥�9h*ŋ8Y�@��~G��t�aRa����G�T'�L�Y��0^�W�����M��3xB����l�>�	���E1`�ֺt.ʾ;}R�� �0;Zܜ��ci��,�N��)��L�R������Ѝ��&���8m �;{�B�V���9��T�<x����]pQ�B�A��/���>Օ�=��d\j���suhL+���.m��C_�C�ƺTP?�5��
��9�7�L)^"�g�z���i�O Z��*��0\V�&-�ܔ�T-��y�q<�*����B�F1�||޷I�a7�^�?d�,�t�?�Q����J೼�B�!��Ƚ��0B�ߊ���l�{DHECo�
M�ěz<��������m
y�'>:Xk���"��a�(�V_v*������/5��:
I"���i<���J�!s����5���9�v�Umi�ϭ������e��:(�#��eJS����{�zˌg\\^(*��!����Dɮ)r"{���u-�kL��[�V� ���S�	�ou�
Y��
,�0�0
�@���>�e���>mjLQm��q��s�5�ږ���FK��xIKQ�BF���#/R�\�u۱����sՑ䩵g<�i4�/Gr�*%��d�P���_��s���e
tmA[YA[���W�l����	'o\�E#꜍_�R=.�a�����H�pPQ>�&ƺ%K�A��|�l�]W6~Q/����
�T����֮AΩN=Q,R�����z��G��F����K%�b�|>�����h���v#������ ����c��A΃:~�����vT���טc�+��5�0^Ď��8D���Ӑ���B���]��]/��#u�P5=O7�%�^�[�E�z4f�����Ic'�#���]�4���th��n�-�z<31����]�%�aWaw��Ĵ���;=�Z�'���u�k\�V�r�`��d�]�h�b+螂Q�,qoj�:�6.�~��e��6��6.K��-?r�:9!Q��ʒ<��9�^���T��ѯ�D0Q)�06�x����˜�����Qo,�4���V�nM��l� T�jTx5į�o��0�9��T�~��g�d�ah�]]H�j�=_k��EM{tV�yN����ߍ���C���ғ�ۊ�F�o�9Ǘ~tb�󦻘E����k'/:���s���L�q�e6�oT��GO�J��YΨ��O�؍�>�f�{2���zkE�̢��Ը2�?�RYڈ�ؿa�je��i�2���[�vH�Ƨ]YWt)*�������[ ��x����(B�/�9r���<�H�O���] ���n]SI�Q�9ɦj��Mr��ѧ�`�u�/F,�kYtqm���{h���i1��T��,���%��f���{㕜�H�����4`�Vf�Z��h����w�/�"��ĩ�������?���;k���.�:ض�8r����@�E�EK�fd*��w�Us���������޶K���8��'�Yh��~�L�<(�$D� �ǆ4��,�r6�������x�(�j�gQS�w|O+�z~��ZB9�z�,�A��w�/�G�Lj�.�g�f��s�W#����~����,d�,�6����U�ψ�xE~�_J�	��"������j�e;�#�р���?O򡛧�_�zҳZ�h3?F��[Yn�^�q��lz��j��y�gZ^g�$�\��̩RC�����@n��*/J�W�u��*�c�+/`׾jr�� [�������|�ᵶo���Rpb�7AEUd�N�
V5�)��4��
[i}�9��ڀ��E�q1�p�?_�k���-�!PI�#t�8&�VG��KI��$�eƞU�j�P�)+�=c�)�ÀТ��1+��X|�a��~�MWL#�aʉ����v�i?�(+K��χo��+�OH�t��x�Mh�>T�<:�%��d�>'B�ފ��X*V�i�0	/�GB�f�;��u~���zb�I-�\�`m�[е%��*'��wb��v�.�<j��e��[RL�:�f����cvrq)%Ei�B�ρ�������g���b/��h1�E{�ˏ���Lk�fiP��&�c�yp�D�Y�x?����WGn$0�~̆���'
�r�B����Nǹ��s��P�)������2���E�#��u��O>���ʷ��!,Q�Y��OqtVZ�������(��:'~H ��\��+�O���u��yƯ�_��K?�)��ZBW��B��@�#p9Gn�C�,I��spz�TzO�م����.g9�%V��9�֏ O-nI�֧�o$g����}js��/P�Ξe4m����3H��@�;u�Vᇑ��Gq<5k9~��*di�\�7���Ȯ�qϪ=�\o��M����*�S�[����4l��慁�Ѣ�8�rn05Ă����r��N����<Bu�����݄}lwt�x���`!�����J�/
_��+��h�D,�1J��O��hGW�`i����>Ū�Ԥ A�h!փ���r,�q����$��: WJ���;��p穠����^�d����CH�I�mZ�JYe��˥� = �8�+��r�yٮ2������$��}�"�L��^���(�9�.�p�e7�F���=�)y *�Cv�9WW��jf+��ˊ#`�<�D㲒yrv�3߶]
k��p��)`�u7�����$� �W歉�����Tt����EY��lZ��Weo"|O���[�5G0%Q��oo�	~g-ǫ\c��m|#�V��&!2ڳ�x�3u�T1Y���L�I�T(k[������Z��1]IȪ3���"�u��4v�8�H5�n����E]�q-���z�%F�@r��p-`�"x�{VH��w$K-�W�b����f�;���x"q��أԟ��tb�/&TP�F(�o�~��n��Ej����4m��df9����郘����H0���65����Ɖ�RY�'�o�N�I��~��*n&�tԡ�Vm��)�����Qvŉ4�/\�����c�ș���p���D�w�2 ��zT4´�U�Cf~*e�-!�F� !��� Ev	�� ���rL�fץ��v_fB]
d���@'��n�u"\gW��,�-w�N�D5FQh��n��m�����P�NĄ�Dv�)��(��r��jo�lQ�H�o�D��+͝˽}��[5���P��"n�_4R��G�S_��S�˓͈�*�i�n�'��Ʃ�;�?7]q%������,)��`Aud��1'̜&�ӆ[��0�ͥ5�I�C�Ugi�S���6@~Ϻ��_NC�۴t�4N��	؞s�$�䁡��Yb16����A�VH�նx[p3h�J#���V�Y�{�S8 E����������S4���7$�,��?p;��o�kmN�W�ڨn��u�.�c��}�h�J��AB��'��D��x�f��PG �-����D�q:�RQh����\m��f���e��]p���_��uaqm��l���0�����K��~�D��G���rGi%���������iv��;���#͸�vST��su�m;�m.k�c��GR�)ٮ<����F3�DX��՜�{2۠��4�%�hC>�qX��Y���bH�I�yS2#�6�4x�=���h|$�[h��oM=ٟ�B���nm�,1��MX*J� �y}^#�����8g���D�0�+��m��auՊ�����{"<͢�mD�0��������9�J�UD��W��T�&�`�H�2Nd��T6�_���g�l2���h��g*i*k]��1�$XBtm^�1�RX�7�,e,���[���w����#x"�\ ���cG�m3Τ��D��p�<��d9�@�$c��V�U[���H�wd�m6� [�3�L6��U��O+�!�26o���,ݻL�#��w`�W��� ����>�O��-��`����l��t0;꒚���+��Fn�nG\PǺ#Bd�@�/���MM��z�Ѕ�^��Y��C�ÿ
N�q��<ői7r�7�t�Qmf�L�����)<�S�a�v��w����G�X,��Dıb0ѳ�^R�Լ�#�zp��"�z�^���#[����N��q6�
��Į��[MV��A�V��e�A�W����B��xxٽ,"��y+s�,��kR�v}c�Kn_���(�Ϸ<��3N��@�����������T?_�e�ym�&o|!����d\��f�P����ܱIQ���в8
r�T��ME����wC�� �V��
���G/D �p�^����8�X�_� Ԗ��Iu�:��E|b�5/��_��4r�jy�뿲�8�T߼�{����@�۫ս�^\(I��E�ݣ��ę��:�؞�5��5���7�Bn�d��g>0k�k*}�'�s�zF�M=dN�	B�y��ǨU��:G��B>4�/���9�+VA�T
�6�w9�rVMz�!�	��� �z�gn̈�U�n�}T/�!6x���K
_���B�>�,(��i�L�A ��U�< h
7��_�o�����A
��f�b�oC�=�f�6N���W�uQ�W_�B��.'�¥�S3��c�Ql��m����ݭg=Izʵ	�;,�k��%Ɛ�P%f1!���yC4Ɛ�M��E�ٖB�I�+m ŔQ�@[*�&.�tdaRwhBZ��"2��a"RO��s�M��X����=�Hc��j�e�ZWځ6��Z��E;f�{�����������͟�=�ŧΡM�ZƓ�9ƷUr��E=��x�SM����Df	�,R�><�2�١s#���O�����fʚRl�9�C׾EQ֖�����ͱ����K[�2w�C#��sr��_�����%;>��|2��h���slf�g[]��]kj���M�!��e�7�j�^Ut�<��G��˱s����d|����¬���\�7����s�LFZ�}v$�V�OS�#�;BVpg9��m�9��q�۲�o~Ip�����b,���	550M����!w�~�/�U�iO�o��g2���T�R�6��[Q�s�%0/��$�Y�އ�Ք#�"�ɳ�+�y�LU���)��g���7#!�ʨ�hT�5��#k���^Q.�\�U(;��S�˯�8�x���r����"��`�8��V��2���;���{I ~�$_	F���Y��-F6���%O[�H^��'KO��'��:$	
���a��KM%
��oO�0D�[711!�v�@Շ{��k��. ��un�}�q�3��a��X��=%5��%�����J��~#7��v�*�n�>�d��唕cjk�I��BADt��y�0�pC���؈CqmT#X�_۲�S߹�´�R蘫�ū��[��R]T/��g&����@�\,�����޺8��2���+}��2��O�8Xr��(�5@jO�� _�	Q��+�ff��A5�wm`i_҄�:sU��l������~�eo�//���*�7Օ.��^�R	��ێq8�ɥ�+N��;�5[�%�aK0�G6������O9�+O ����uR�m��0�.�w�H��!�3�W��RsH�U��Ȕ������khނ[�tI�N�(����	��b{rj�t��T��h���`v_���Dr�m��3�ޛ~�;_Re�����t��������cIN���R�l� �Tj5#a���o�ː� �X������-L�yMՋ��D�'��V])�x�ҿ�]�xd�s���q��쐠���7��^���Ƙ�0|꼱��Pb�G�#�������% r�|�����텇Z��e-���L�ǳ�s2���C����kO�7W�Js��G��6>�2X��W	mi�f���@�Oh��I��҆���Ut_�U�;��*�q�p� $r�D��߫�E�BB�Ύ,��I"|���CP�$�6~�ѾP���G>�B��~`~�WKʿ'��Iڪ�9h#�}��#i�����s&�7@q���0my�&��,�/J��a��T��^+��o˩D��������V Y�G��6c�{4|�%!5h��Ǒv�]ھ\��H�WX�=�����
5�j�F��mb�AMY��x��K��������4S��+�@���BR�W��s8��_N�`��ZV3{�Zկ0��
$.�%���p��� T)C]�A���v���Q2#��y���f��r��$)4������Jw(5mCbc���D �??4�������������q3Od.��J� ��h9I���ة�_�KVN����H���s2�&��k�9S9ɍ�X�!�:��E7{�u��Ӻm'7щ�6������]"����w�$(�n�9ڃ����'��
��а7��ѿ������P	��y�y��	[\�U�_�:��ʎ��7�0U:�.��FԙLĢ����G���<��e���^�ME�y�^����0�jf��Kc˓��N���� I�J�]7����a3�٤l+��}XO�;�#�m��W�����
Wg�*=;v/�@�<gA��1u[�M��ⷌ��<�:�7ф��F�~�7Vy�'N�̥��Pѽpqlv�k����֩�-F�X@��W��{�HCp�+���=���^�8�5Q�O�.e=-�[�y��D�A�q�ʫ�C��{noGj���$��j��sd]) VY���} N^]l�8�)�\��٣��]|��`�L���}��g�o��re (�s	�d�<?�U��?��S� �a������&���#eK���E��:Яm�l��hp��9�S -3�/B�?�x�W]�e'DjxO�;��vͽKKȄ�=����1n%��C�z��M���-gV[�\X�f`�QGF�� ���)�ٔ{�q��ƺm�':W&��<���FK�b'Wi��I���tie�|����K^��ôe%�~�g�O��v��/*�&e�rE-L��-�B�+����6��/Q����m{�F���`bA��*w�Aߐl rI����F��p�2h���>2������k�1����8��26���r�Z��-��gkBX	slS����(�e�R�Z����x�W�3��	��Z���͆�;�0�u�U�9�>rK#ې��i��)�o�:H:9����9�f�∾e�;�ч����o��}�霯�(�c�C�� �� xC��y!������-~��5�}t��f�c>�&ׅLQ����`�N�E���1Ih����x��ք-������I�:���ĝ�H�Nr3o��&]��v�R�i`S�GQ�sR}$:z��.�U� U����,烄�����R=k��F����w��κ�:'	2eF3�2���t�p�"��M��(=#��Y!��He�C����e�G=�*�3E��t���_��,�T'a3���`Y#&i����H@�$��`��("���b����?�c�
�R�� 7�bƷ�'$�w>�h='8Fo���D�uS�ON+w*ٸJ��zmC*�-)���՗;�i��R5&ã2>���V&�h� 't�8�3ݏJ�Z���=�i
��%��|2���
�B��lB��R	hNYd\�J�S�H4�3�����CD9/�k���H[I�No�5c��e�]��>��o'��Z0}�H14,���S �6���Fq�w*���|y��<�u�Mx�'EtM�Xy���]̑F�tP%�?���1���"���[���}����c�����?q9kkP#_�)/i��͸=�X�0vu�&0sN'�Qfi� �]�ql�"]Bq	�#�d��eH�坁�������4�>�-�8��#�5-��/�\��N��!�4C�'��t$�h		��)�:hI��S�&�NDH������,a�-IM��Tg�����͓���Bم<�������ՊM��b��z����t���N
�p��$J{#��Y��� J�A�Ar�Z��|(܀E���OK��0,�E��k��J4�s��@O�C�7JI0&�~Y�+��	�d�̈�Jg��,�SI�\I:�m�i<pA=0}f(�����L��7�ax��vPA%w�A��nwz]�lR�yEcpC��Y���:b�sWWLB���n���W�g��%pY�$#��2�I݂�q�*���*�:	7��!�Bc���+m��;<H�o����&�+�	�5`�O�	�6F��P�E�Z��_Feg�ɥ֞$Q����$������ ���긖~��;�A��g�IO���j��T�啢�ЕJ���?Bi�������s���YhMPe3��I���+,�2k��Qf#v
i����}�<$��
� ������7�]�a�E�DD�oς@Τ^���\�,B���|�2����}W��)3���a=[I��*���n�@����+�[p�*�٘���
�����(.~��)�@p!ܛhiΈ�Vlߎ�LjH�1Lo%(�f��"�ު����ɟ���G%��󅴌(%�w�N�o��K�2��~��n+A���:���x0�#���Ӆ�E�a��=��#�6"�j�c���;G{I��,�ROib�Y��M~����	x����x�C�}.�	Ba�a
!�t�AW���^�p	�XNU�;Pzf���i�n��T���	�X*�`s�5����Etm��=ǩ�`{����qB�IJ�+�`Fѧ�`	���	4�yU/� �e���̽���L
�4&��AE��LQ_UyB�[��KO�C/�ށ��VsऄZ۰S>_�-b֏��ʯ
0pC�@y�k�ا٣z�*�-�T���}|���\E`�D�[Z��6s�Z�u�⫀Oi��~�4��ׯO�ބ�d
��T��U?�a t�d>�z�W�",F�ҫMd�t�*�K�<d.}����j}{E�4w�Q���&���/�����	>����*�Mb�T)�]C�H跢�g���j�Ϩ����K�韰]214���Fo  Q%��� �u��x>{y���AeGy���<�*Ч��]��L�|���m� >�v,�Щ�0��A�205?S���FЃ�5�~3#��t
'�r�}�Z�>�����v)��&� ���H�ą�5���)]���$r(��ߔ�ΠEꊝc�q��Ѯ�L���M����M�l�y��
��/gv��\Jm�_ I���f��#R�����@7�~a��N�3f�Mm����I=M�`71Y�H46w�(�����^օ�
�8A�3WN�D���RF\�dgz� ��d�7���C$��s������T����%�}RA`
��vOf�I��z��\��Su�%V����F�O�g'{�T*AZp��p�����H���V&���6CF6�me� ��MwVa�d�� �@
��2c��Ov���V|�nT�4]��Z%
�$�/�\sP�5h�h_�R�t~ wܫ�i��[a�6ݘ0۪��׷?w��x�;���� s�[�ʂ�8�#�|��Q([k��N`��,j�P͚�Uԛ~�,)�V��0j��Iԁ�mk�>�X��ŷS���E�90�o����o J�i�P�1����p"����Ar��؆�D��sq��+�l�5��^G��uUw�!��xq�����i2�t+ʪ�*�L��휘}沱�����!�&kkI)�m���x�T��m]$�Ӕ:�L+��^mJi�0����k_���-vHԬ\���˘�e{��/���@�F���0�
�AҮe�pCO?�bEw�镹N�K�c�T(�w��d$�Y����g<��#>�bZ\�Duqe'lQC�z���Ʃ$*�t���*X�oã�~U�!��*��ST��i>�j�!	M�~-g�R(�� ��.�)�Z�_Q�δ�7gQ�-��L�|2ey�#�b��I��)�d���Y�U� �����q*�����A@��?�n��e�x��I���Ib�itT���Rу�;E%jn�PB��Rn���s��u_ ��a�ܮ?��4OpF�/ӵJ
�rm�3,��rJ��Vd�`v��ǵԥ6&p�b��n�©�#��}�����ۃ= +-�Yƭi )G���M�e����Ր]@=��g�k�;T�@ �l�Z���o6�)��e�%hG!SV��\Sj˽�a�6j(k]Pϕ��?&W>��˙���VS?��}���Кvi��~�aDd��L��]�7���)��dd.{+O\���SW�b��iEs�E��E�w��]��x���mҸ꣄��1�R3>8�����U����t���s�U�w�;q=e�Ẓ��n4WVsܗ�$x\)�񐷋����OB~T�W`wuƶ��k�sD��,
?�S�Q��{ܴ<���yLJȩ�����0Q���p�7�ޘ$�UG��o=p,:gA3��&�NS�o����w륏���b��!6�u���ճ?����9�	9!�b��4qI
��,O�Č��°��H�"\��4ut�ʺǥ�A�`~�I���̹4q�S�"`"T��=�(�y䴚B1���|?�
[
�
_���`V�M�;��2��4�w.���WJ:MJ�#�XUk�a��NM����ߩ)��ږ����`_�R�4�=)}=���P�GT<֨����p*�'-s��R�R]�s��U��J0�śbi]l认��{m,�f�d����D���9z*�]�)�?JIC��M��c%���9��<Cx� "$�s���/�:��|�0;�$���A �b�W��$&�<6>��~`�1U�.��
x�(�v�;t�g�6_���Z�;�z�1�^�����;�;J­���K��!>�j��ͽ��] ��U�!9��_A%7q��e�����hy���؅�$�T�#3�=�U�7_B�̑��z|�[
��ϯm�3�c�0k/��o��s��Ԯ���-����{�(TX�Ȳ����o�d�s�;}���>������٘����@6���e{%�eA畽���ׇ�K���~�ǟ�
������58��Q,���q���TU���v����0�����m���utv����5�mC�N��	�5`�]�©�1����Z�BR��2��I2�Qeu��n�Qa�'m�-\;�-��
�-�s�(�]�6�˒��4�9ҋ��:INp��͖_y�f�����&ɐ]F?߾�SF� ��^SL��X�Ty�x��-#���oC���?a�c� ��o��{�>}��+dOR�8���i[�z�W�7g��:� �c�������T/΅mD
<I���5���ൠ��+�ʒ���=���/]L9�yb�����Ty�󻙺|>�����!�����&{x2��g��7�̶����Y�<��ۭ��7G�(Ѱ������,w�/`5��6xC�I|��,D�S_�ç�L	S�$X;��\�Uv�usVC���L^>7����8bR���!�':&��"���J?��å�*��k�4��J6`�5x�H�R�w߃'����Y�I��Q�@���Y�K=vi�]��e�$�#@��������,�YF�vf܏�;����d�_�� 德���
��W�NK�,��Yt������U��<�'�h��>3��U�u;Z�T�6>�!i����s��X�$?FSb�<��m�T�C\Ry9����;K1��w��3��t몓�1��a"p���-�%q�݃�(�AB����W|/���U$U��g�6At�H*�~��z���c������4ڏ%^����Ԧ�Ӯ���j��H���@����W�q64���z���Q�!5 �L�u�`GT���ꏶ#�ʜ/D��b#( ��6���W���v�J�a�y��w�|F�U""���
ɳPR�(J���&�޲��J�x'-g_Q(R���W͊�_���x�F��ւb���\���y��R03*���n=7���h�\}2T�������2���}���Ȯ���wÌ2 �j
��KT��<Z����xc��T� �
.�X��T�v���b�4m�kR����46wQ�4�����Z!�}��Ȉ���V��Qz�v��M5�E�5��Ҩ7�/]��ĵ��.�.>����`�7��'J���k�brF��F�x�=w��i��R%p�[�J�Y���G��]?���C�b�䑍�Q�quU�Z��������A2�� �{(�����V��4��K�J�$�� ��1�Ӹ\0g�1��v�����ahrW^�DWTD���O�V@��[��y��
�YQ���oJl#XPG���=`���R'0�|�9_X�f��*�2�{����Z�']��a D�Hkr�;��-��\�;g;�c.���'���Z�b��D�d'~����ZEh���?�x~Y�����K�N�2V�2�tu����ɹ��Y�*8�K��BkWs���#R�����2�a����;�J�9A|��܊��x�ד���7�Ah^JEz�ik��>\�x�>U[��&�Y�4QE����I-�׷-��~:T���jx��-�5�|����Z�ǌ6M����-_ʨ�O�e�$1*�	�=d�e3$�jk��챦��4>z�ɧN�,����h"�r.Z��V��P�\ �0u�|��{T�k`��t��6�᏾6�j3��L��k5m�^�x ���l1���SV���!����GN������0�S��(g�?d�����~qՅ�<��.�V�0���#�cL}��&�o�z2��iDKׯ"�O9�#��d��\@ �����n�5��z�#<6L(�`�?�|��:�l�%w1�_����Z4?0́'�8B��Iq���P�Rl�{�/�8��d~oo�a#W�O�I>ǰTߌ:�Tط#�h|a�ҋ��T _�2PB7���ˬz����`�!��6\���A%���2Y�Q����!�5�ɳV���f��p�6}<RR=���F-z���2^�\;I@�;����s=���wx�#`7�����~Ĥ�&�p^�N�;�6*����S
W���+	�������V��D�NF���x�[!�9!\|@A؄�-KL�!HK��g���'�d�16�Uo3�	#"3G -yx��_��-�볾�%��Q!o�r�9lJ/��7�u���܅�⃖��[&�r%󜯶����(?q��yz5 |�>���&b�|����L�k�ٝ�A�����HI��	t�Gh�\�VINc$r� ��*�"�.��>�������!��:�:ӵRI�[�gr��m;^��:	&���nb�[��ٮ���5����~ }��$��n��(��� ��`~I�ɼN*d�X�pı�%��v���mL[�I4(��0Ή���$�2����;R7$b3;F���QKJ*��-;����<�/-��f]r��=��K�T�j�RRB3V��KC�#�]?89F����h�S<�-8O�-�	�`�?_��
4���Ǵ���@� h�ƴ)�"0w���kL-��DBc����_��S����A��$2p%�آ�������\��*L�'R,s��i{���ĭ�Lܻ�7�2ݭ����Z����f�>�6��ژ:�޶A!�-��ѝ�v�������ӗm=�H�ad �9�(���0m'Y�i��U��\��L|���._9���Ne�MD̾m�]/
Io�Y�L%Q��R9��s�A�q2,ۃ�����0��4�ir��������!x��`�IiG|mG����OV�*�s/��`핚2ew9�W�f^���Qʪv�J�8��5)H�{W�۟B��sw��]zL�AЗn�p�o�b9�D�V��dbhۙ��L�)&w����>usž*��+t}ټJ=�I�8/88
����-&�!�8J��s��Ei�;g8 �欉Ud!]p;�������vs��0�2R���E�K<�ہ�����u�G<̐�sH�d��FW���Q���Œ%#f~;PY^a�ɐ���e�5��}�s�\��7e?���y�fw�۴��{�B�d�}�:������ �+�ݹH��3�M�oxa���KI�V��R������G�^��_Ń�ͫsI.�~�l���d�`7~��(.��ɤ>q����9?��4H6�¨��{I�#P�Jf	Ub8���T���r<��F@ĥ�y7{d�9����NP'(�\�¥�z{��P�<B��0�A�z���Ss�"�m��|�ypI�o���-{�\������و�,���m��aA7��h��'�:��D=���XZBxt����!�5Aޮ�=+Q�����JU�j�Qz��ޛ�o1!(s�}����XEz,v�-���{��}����ė;;BQ��9[b�@���E���.�o��W�3B�6�!�7�"�sȇ������o!e��gh���򗞥�[O�,|���A��U��:����E���wG�$$W;�������xD�Dx��{�%��k��i$V�=vD;���ݨ����>��&��=1�>G�<�/�SMu]_����K� ��O�_�8tN�gߘ�i�o0yg��[��Cp�����E�:�������0��)j�I���Q��x��ޓ �j�ϡ�P}�z���|�&;	q��v<�@�����#7�f�7oL���Ť#jN�!HlG�%����<��ʘ�[����(�3q���z����,7K�]FD�1���[���N���[���\.@�Yd�G�g
��'g��x�����>T��#���e��3��}*�HP[sɸp�t�;���2���bk��ǡ"���)�N^����:��J�P2q�Q���G�
��y�����b��;��0���v��fK���\օG{;�-`xR@�_p�y�l��I�<{ߵ�<S����c�h�����]��0�,��u��wNב5B�1?!+�t?��1e:�Bn�_X,�E�c[Sk����ј�����_)I2��wM�8N>�M��)2���=��D�Y��!?�e���	ʅOB��m�H���ԠZ.f���v�d���E�1�� C%�h���3��
R5.~|$�Y8�F�O��z	q?A^B�/��q��ϔI�d�_+�"]�����I�d`�&Z"���z�ə]�}�PXe�ⴺ�Pz��2�g�v�y��������8�Kw����3*����H�N��>'s����R`����(���^%C*�@������'���q�W\~7�~��!Ε7�w�R�d�y��S��::��x��/Q��/N<��H��̬�Op�2�G�1�Mv�䅉�ᭆ�����'�9d�F�tC�5�e�O��t���sZ42x_>Sr��B�o���&m��qt�u��n���ipf	�w*�m��.�����@���u�&-L��xAB�5WY[8�z��l+��F��A�Gق_�"�h�^g΁�p�򜞷wQ�<F�`r�t���|�%��2�y�MF	�2Qܧ��4a�E����L���lA���&�R�m5�"P��`�^�#�tm�cL��z�'Ճ`�n�������3����rA׍
���#�� ����c����%q�=1|#�h/�h�w+�eS�*�U�{wBɒ2g*2@`�1�o��g�9�?H���!z��&Y�{��Yp/  D�'��-�</��)E�i\�PA�Oo�]U����H�m5�4�I�]rY�ܱ�s���|���i��r������!���!�a��a�4�\;#ɖ����b����C4t���0},l�nG&�ڃ���R�
T��̯�S���Հ4F\�iH���7��0�Ǥ�ٌ�:�� ��
�ޕP��ɕ5I.�,:�bT�$6���E�lʫH.��44M�?�c4��O+�$��z�ƝL^�Y�6�
�3;G�BC>�����X���oz���5j�{��bQ�젰��JBd�jF@UM�^�I_t���1��>5�m�|C�Nm.�O㢉������ �<^��p��H�j�(�<����%o�U5��ta��P����DU�g#KE���<\���d{ɘq�"�UwV�����*l���������x<���F=%3��n1"���#�A��������P'�b-@�L+=��pS�0�[����o7F���E����h7��d~p]R��4\��<����ry��-����i�ԋKu?Z-�O��V~pu��������$ոĪXh_�c(��>�K�*s'��sz9�N3��z3����`q��Ϡ���~$������OP�(V�A/G�v��W
�j,�+T��\uR>��ż5�XR�>���8I8�[�-FVr�˦�U�Nw����"�
x��)�?҆8z����!�ȉS�W��O:^�BӒc�w�@.���]�J�,�a�7 �sZQ� v�t;�b¼���kAR"*�?�j����|g���
�Ȏ5�Y��`�)1��"�ĝ�@���8�Vu���SQ������^޴��gz+��+T��e��R`ޕ|��؈��,����/���h�3v�<�C�����lXN@{r���S�q��Sn�ݑ��	1&���~��"G�^0��i~�ii���7��M=Yx6�)"��
�Ou�r�+�:=���
��k^�!+�п�J,ǭ�և�O]�# R:�~����
�c�$��S��5��:[���hC�χ5p:ml�� �zb�?X2�5=k�O����J���[h��]�g�˧%OV��7'
�Λ�b[����O���~��oEOd�2�C������}���ܕ,�n2�,n�@>E�AF(���77��<+}�_�Z!L���Zd
&�4#�ѬA���U�e�N���Y��!�-�Ek��ȀP*�Ҭ���1r��{��B�|��h~7���<�n:�-aʦ���֫WV����*1�POD��ö�5�<�)dk�`ւ�޳*���+�I��U9�����1�B�(e𡩣�x $DSu�@�B��ҍ��_�Rx���4�wi��mT!���.��E��r���D�}иh	�՛�B���tH&��$$��V�T�9G�(�s$��� <+����S]aQ��<��ĜD��Y��b8ɻH�M��Ǿ�ӹ+�!�Ab!�PՒ?U��8QW��-T�Y�(���7h;��mF���m�/m���ë���YK�zBŠ�t+(���^xbM�7lgXn��gi�"�DL�Bj��j_��W)���0�=��Pvr+�z�#��0H ����H�������!(�:)@G�{v�
V�S��{��y�f|�j��t�[DY�
H1��������.G��}s��T�����5�[��k����^��������h[4�Q�vC��ՓS2'����X�E$`�I���G���N�mύ��8.���ݱ�
�0_m%������l�w�j�d;���d�;�4v��w�C�]-xP�Vo�|�������:7JEO0�+��`=6�i�9�JVc�4K�'I�:\�c���,�u땋�[)�7UQ�����BM]SR�H���|q>R�*��|��[-�EX�
��9J���l��id����b���M�e27�o���9�LZw�[C��=[���J"�Km?K�4��h��&&�rl���U[�DZ0�p��S��W�W�Ry�+[vd����K����|��NmyU��eB��И5��,��������_1O ���8�Q�DʷeM!�;�r��շ����Ӛ�i/�G�Pm�ÀG�D��b�pe�#�^'��/�-�p�3՞-dv��I�h]t09ܞ�����0E�S�Oc��5/�T�=/��ԯ�N��`d�a*6�T�����>�T�`��	Eо����8ƏP.-���O:B���$&:�
ƚH�h$��[���I��y���1\.@���+�juj?�LcPV:y�0��(t�ߋ�Z3%�-�5��9��L��x(�Úe����g��0��Є��N����_)ڥcȵ5 &���=�՚��A�#ue���ɾ�����!f�J�]������w��2&�}�k����q��5�E�PE�"`Ȍ���Ѫu���<N˼4��������d���
J#�<�1�H����+.�{N�%F�Usc)	�ߞz���|�~�eT�Z,�Oc�7}\��*{%�;/-��%�JG����(%�`|xtu�}���S�zl�=�,,��Z�A ���:v�i�-;�+�
rF�P:+�M����9�������sϧ��4�Q6�����><iD.����~y�h!�p���lr4�0��r�!�̅63p$�ţ�����S�+&H<����d����k���;i��~�2j$UY��/Π)���28[�VS����[�+h;]�0rΙ5�If��1�i$9�v��n}�p��1żP��w3����:��������56��y��.^I:�R0vt��l�BӍ܁t��Y!`&j����(]y��{]tYĮJc�+��0ٿ�R��~ )�|��5EW6��w���
`aHc���������2@s�)SjꥈX#����F�s��m#��qA�aBP%��2Ӛ�DR��=��i�2�4Y�,�Q��e��b��I}��=����oam=��x�K5 	��K�E�[���EŰ�@z�e9s\����H ^�ӄ���~���W�����#��v��ĵo�Ь�q�D�);�H�QX,����͈P��2R�V���sp
������8���#�L�5;=�z�hm�Sj�y��O���8��<zs�&ZP�����e���`.p��-r�A���x���g:�����C3o�	��K�����Nz7?L�袳���c�KTw��o'��8�8i�UZJ��"�ɏ��O�K���I��U��ibz����m�4*��3{Wq�I4 �h5�Tf�d�<s��멵}"�ngD��}��2h2�7f8��Vn��B��]������{c�%J�U�J�x���ck�S�X�t����#��r���f�7�qR���_#ˢ����+��@xۦU�-���eO�%RA}���a/w�BF���w��?j_0�o���f��ʠo�����V�*|ՠ�������/4OU�s{�2�����9�����ޖ4�w�-R�f)o�k7/�Y�ys�Hh���S��صH���yR@�묽������u������A{�;㭱�;�I����v��nΏI�V��V�|0����UGd]�?���V���C����5��yz�=�Eme��0�GRC�!2�Z�u@"	m�1�x��|�Ec��|�?�Jilf�?�-,��W(W��<�`P�3����- ����������볒�Ryz��B�[4�K1p<ϝ����%�LI0���ٗ8�ϟ�i _1IS7��L��4�	iu)k���"�6��,ʴ�6����x���EЭ2»�x�$���wf嵨���中OO��4hK�RB~�
��l	��kg�}J\�����*[�j�P��uˌ�r��*.s���|���e%B����N�A�[>ŲRV#7v��X�@��t�딥!`��ެ����|!�ߝI2l ��i�j��=��h߅�4O0��Lm�o[,Ћ��F�?��lKa1��?YX��FG��,\�vL/�gu4\2|h#.��f����������2?�b7_���I�ZM~��\f8&�a���W/��X](c�۬�x�e�V��0o6���@�-�<L[W(�[�����'	>X�L;�g��Al�{n���U��C9��b���g���`�y�T�aTm,�� ���l��ח��0CO�<u��\��S��Yrg��޴WW��w�W�u?���P�<�7h7����p=��>F���*�o9�� �#=&EV8������+�T��/��f%�M��]��f�0�OK�Uo=�.��>׺�a���8��T�`ؗP�z�@�E���RpoK�)����3հ���4�	�$��ro��`��x��7LF$�L�7��&�:RX�r��<+�$:���u�m�|��3:R9�D	��L�^���z=Mx*���C:�n(��������u���MW�=���Q|����YyCK���QO^�����8�EP�1J�0D�"@|<5�K�K�����]W��APt=P��;��N@l�O����K,��,Q>�籆ϧ���e�|�9ߧ�����,��
�	Z��Z��M�`g�cD���)���Ȱ���3��X%yȱ�ҩ I�4�nJ����_ u��/ۃ�8���{]d�A��%�~1��$J���	!���A!�����Wّ�k$0کU�*A���wpN��eu��/�X�:s�*���B��)�,ԟI����)DV8ڮ��X����ghlZ��O�y�O~T>ZL2����8˶#�W�7���7��2�5��������H�h�,V�(D-Wv��R�t���"s=�>#����4&zi�{��]\h�[8���ǵ?����]�hi
q+�,О�LI	�,,�oT2
������zyP~e�|;"-[�����=�ہQt����9���3�A��a�z��k�b�\0=]	�UAr�
�|��ר$I�����Lr�E���y�v.��r��D���ek�uSb��~��4�%��6?)� <B�Ç�Y��Ӈ�cU�a	:���@��vs���B �W��������B�}^+*)�}��L�#�1�^gxSbz����+A������L���r�y@T�9��+��s��%��'�R7��h��;�G�jO������l�(�;7�a�ѧgi�9�d�c����^&�m;ȈjeZw="bP��Kk�i�"<7&��ݰ�B��?O>f�mb�v�>�աP�I��s�jodJ�$��5b���9��Up�DeƯ9�6n��wO"Q�;�ص�zZ(��iF�q��vO�l�0�ǒz�#;0'ܤT�)��x�5�C�ǔ�K�2[�l����@\�;f�V��]p�-*,�j[�n�@��W�fF�)RvJRp���=l���A��d�Q�@b�q �PtPkr�����:_e��=���'2d�xf�ؓ�Uҹ>9���|#���U&�a�PAc��Z�E���oHg�����5���=��(��#�����lH/��${+Z?�2녑R M�OwAsj��5�9��+�O��������z�z���C\Ȯ��2G�nb9�~�&��M9������� :ϓڏ �b�x�dgƏ���뮾�P/4Wq���k���@��J�)�>�7"�p�=Ь~?������z�Js5h�c���#��!���� �w7�<�Y��c�{���C��)�j��� �V��B��|w������G�p�{�P����H���i��A˫C?j�ZC�,N��wv���&V�����l�X+$i��AF�G2q���R�^%\Wݼ�5��|�� ��1^|1���U�濆*��u��q��Y'C�Q���|S����)5�xf���3;s �>�_�=Z/�^�@#b�JZ�<?bA��s)}H��jt)�*�}��RI�oG����r(�A,�$}���Un���<�q+o�4�K��I�<�mE-S�_��|bO���]B��x�FMD�<�~����6��`�i���6Z�u��sfg 'ظ�ne�=,�w��? v���d^|ue1У��S@~�X�6�=�:DO�OVH��[�垪z�����J�L���R�sb�c���0RR����DrY�x�ਯ'
=�&�v����ٿÜ��0 }v#�̈����;��N�*^me��9*��DG�t���ʡ�V/
���j������A��*p߫�RC̨��=�7�ώ�/��#�c��o�A�{( 2�q�<`"��P�v�����8t�}V��ųU��*<���C�3G����O#ں �^�$����>6��a�=��(If2BJ Ŏ���>-M��p�Y�韄0=QBolC�*Hn�o�������Ĳ˰��%U�Ӳ�m&���0I�7��9ԹF�r��=�?��/W?�PP<� �X<A)��4�F{kT�[u���7�٣��L�̫5,�fD��n�{R��x��%U�U�������б��~ f=_}�&��s�4~���)�T�D�z�����(L9m�PθE���\�	��)"�P�L7��z���a���kd�o,��避�ra�<�a�nO�!��Ϯ�sA 3LU�A
=WoG��3�k�Xz�j�?=�}�ｬ�,3�w��4>�"-T��󛿴t�#�|�R&iR��R�t~E+I���W�)���+�Td�<��� �N	�]�v�`"�Ω�FG\E�2�e���}�'5#%�]��^��(�RY}��{�V��z���X,jQO�5�i�Y'N\����+!�?GL˓Fu������%��(�ϝefjN[^�"�v��}*��j#;����!�(�`�o�s�u8(��$�{6��G���f!�ǘ�.��D��,�%+i���k���՞���b����Sk��q&��<1�%��z����!X>��>�F%jm��ϚX� F+޼����ю��V�[����(*�I4�/�>ЕT1�������<���,��V�d��v��:S!�� �>��ܽ>j�^��5��/Y�g);12IT�옭���Gj�-��m�:��X��G��d_-�a3�x"�H$i�U�!��c��4�mVq�k�|D��&$*\�1������F>jQ*g5�鑚��nJ]��;�hqR�Y�9yT;φ Pd0�;+���wU|7I�U��5?-끳�9�mTx����T�XZ��@K�!V3�FV�F��S��=	1߱{���G���î/�F�`~�m�{�����t�j���l�U0�%gW�)'�I���FO�<�u ��̡̫X{�;�ÌC#޹:���(�q�桸�"_f��:r9#w'�1?ѭ��?1y��jrG�+�!W����������2����Y:M�0�?�"`&N�c(��I��̱�}��]��)�`�`���l~Iw��CC�v����ӏ�=:&A�1���
R)����2�������[t�j��8����5���9��m�7Δ�֓��A���ø����<�\�1"��M x)E�[�+��]��@��ɯ��h���y3A�:8��7����G������*�s�YE����&�2y
fo��]���zP�")\Q1�â���2�~[��]xȄ�����G����\��D�q�!Ι�k^'�����U9��	F?��i[t?$RK��x?㘧�<Y�[JA���y݌��t�I��J�Ƿ]�6QA�%��=��Ab��������;l~�Lx�,���g'���9�S����#�_J����5� H)�}�b��g���?�_�
ŀ\�����K���Q��R�%��l}m�%�䛴�gtx�담�ڲx��Z1�����w3P�����|�54pl����}����-�[Tס5�!X���M~S��Q����nK.�84C�o�^��a���<o���в�0z:�Y�b��!.�kEo���j������aYkF!5IjL�z
[S����Md7CkT	ly��j����w�#l�҉$NN֞��G���z���i�Z�:���K�k�c����� #S��"cdm�l�E�5��b�J�x�$�a�w8�#�QZ�rHj��6,j���kh����
�D����u��*|}��LjH��t�.x��d'?0�?ktc�,�����ES��.�V���x�[��S2g4
A.�d��u�&�J-�`ӈ��ec���E�J��K��	/¸uc�c &��_��!ɔd�"ʗ�E��vH-�IF���M�k��r���7Pp�cd��XW�|BQ�j�<��H�D�]��i��wV�=���[I�Nl���fI��{.�INscl.n}�6����V�P�C�Pa���?�q���!��%
��M�[�t��w���tVe~��W^��Y���pU����B�p���d(��������;�OB�����BC�Y+p6�O��A�o�#�*���#�'�L����Y꫅��k�?�rЯ�SD{
2�(�4�W�-�"���(�Nc^�~����a͟ >[.��2��)l�+Z�X��8z>/k(�f��B
Ɍ���Z����8�����!�FGari [s�l�AM� ������Be�)�D�,��!�4^�I�yT�/�Y���_�	��o�䴅�: �����cCS��ں���y��wj}�PKR��eB��B��:��a�]��;���4<j��P�}/�A'&�Q�E�$(�%P��J�7�0_�F�K�'��2�{�L#L�^�o�]��)F�6*���A�g��?M^-�r�w_�0�жKФ
K,bȽu7-l,𔤦�0�WL9ǁ�G�]ov���$���C���3f��G��t�,"�Ӊ��:E�05Db�j�D�_ʜѤIWuR���kU�S̃O��+��j��2�'��dL�=����Q^%��k�<<-�CX�B6�V�̝�⿮��w�)����4��$�(�F�����]28�T����"��"z9tKRԵ�������p���~L��ib�4���D�w{��
ODL�h魧X��9'��i�n�@�����pE�R�)��s�i�u����Af@�V���������`�\64�f(fai�`t���Qy�(��w��%��8���Y��
C!v��5�Ջ�G��������9\����0V�J����z�Ib��%���t��&�BZ����2&�F���g�6g���2D����`�����v)2�:>C/��Q�l��ȓAd �r��+��I�Ӣ�����P¢���&
0���u"�Ү`:��r3�|ko'�����3����� /D7��)� 1X�����۷�1h�����v�]5�����&Ŵ<�� =�1c��������G��� 2���8t2M�4�����O�z7_Uo���1��E�?�G�B�'�	�znq樂~4aXW���j�c;BfsO5I��L>J�9��X�r��D|�a�!Ӣ�t��xkP	���fć�f����r�F[�I��@�X�l��;�Wf�t�8��+�2��4���*%B�ˤ<T_���Z��;���g޵�O��9sK���-cl?f�'R�a����]uZ�Q�����S��,h]��H�6���gQ>D�.�tT%$�����|\s���cI��sy�H���oق	�Ց�nq<كh���p�s�INÊ[9"�:�d�����.�:I@�MH��O3���eh\)z��?Ӳ@�y�nR�fd��f� ��>b�
"e�R��_�Xn�koƪ�@vĴ��.��e~<�� D��8�I�5+���-��ʤ.�DE�.u��������F0�H��� XFF���^���;E�>�nmô������~Y6P$�lxo@tW�i�do���n�u�ڣ�T��:�����v0�_MZ���T���H���$E.eI^��D�v�	 �����o�1�X��Ґ�n��?K�[�y.=֟�f$I5�HZ�7�&Jo����5%%��Hl���z���T���d����Q5�W�F��u2o���)p�u���{N%�ᠯg�:E����,�ya%6Y�#Nv���˻�85X�)^!��P�zD$ʫ�8�����8R�+a/��}�+ȕI���M�L��*����E�#n(���ڲ��uP6�K	��e�U(�{��F:������teG�6�OM�#����.W�Yd���юg���S�;���������CbPN��F��Y����|*�&r��uRqO��{u~׿tU�)�`��]"J�t	۵r���b������M�^�f����Yv�yO!�I�wN���į�|1�D��[~?���f����ܟ���7�C� ӧ��t�ߏ����,I���+̤߶[��t�����Q�=�\p헰K��'�U�mU�κZ�����CMrMb��L�PhZ�]	�|��X	"v�7��)k��;��1
*�̤�Xq��G�a����5�Z\��E���G���(%���f��*5��4X�Nʸ&Nk�js���Ը��=�ٕlG��u���}.>*�W!=W�Tw��$K�h���8�A	�E�e��~�%�qx���R>M��U������uϳM8����Q��U��E) ���N� �χ��V�ɛ%��c]C�3����.c�q���[����еMVП�Y[O}�&\�A�)�wf�r��l�������ɔ9��VT��k�fbF�J6|��Wo�}l�.���u�����$ץ�>�|��l���<W#K��t�{DШ~�(1��e4$S,&�.i�q<֛(��M��&���a��e��,�2�!:GB`F��t�
�G���8�"�M-�s>7�[�t9�e0��)�qv���M�wm�d>���t�r��c9��xr5��v�H�����i��x7dw�g��4�S�i�d��]��#X���[n�o�t{��r3���z��ufz�6Kl���@M����=K$
H�7H8$J9LR��ߙ���X���<�膤�~�7o��b+�)�C�&�,e��,� J$L�\'���C� Q�ڿ��W:�J-�?k=9�4�"Jx%���FY�����ߙ�b�����E��d'z�åe'5V`�[Q�f�����%/��~P�e{0&?��E�wϧ��YY�$�G3"|A��F���c����l�%�[r����.ư�(���NTvt�b
���2n��xA�yC�h�|E���3.���q9��� Rs԰R���{���O�]� ��WX`�:��}3�����%_c��ZHw�L�a�/��M���^R4K��t�<��V��j�Ԣ8��B3�.�C��UR���i�`���9æ���:	���{?�[F�b��Í���)�:0'k��I��2�Ҳ�_���>�0��Et��1 ��O��)XKaҍ�u(�n����� ݻ��h�Xa_�6�rR���n����}���?Ywh���45��k���EV���8\OKf��9J���]���!Y��%m"�h{~?��(��
��� e{P���|c+�P�Z����xb�]��y֊�z�9L�1cC��IL@T�?`h4�Thn�?q��4�$�k%+�����U��� ���XRk����m�05͆ڨ7qpj�G@��eׂ鐪�}d� Plh95�ϕ�3��w<����|k��b�iXb��Ptf�#_	�{�7��dXr�����#x�ODDW,�NP��{voj����YF�)�v�Y�>�����f�[�!"@�@1Y�O��*+j'5=Q�z������Nt��O������S;71�guv4�) p3�e7Mvv�[��N���N8�b��?mQ��Q�p(A���/ \2��n�<z���.�������w��C�����A#PM�h�>��>[�G[P����f�I�w�t)���<yN�<��GB5_9�G��������v�]o-��� И�j*�.��t�����5đ��^���x������D�gنmH�LӱX�NpCK�/Kx���L�\b�&]Lv��пq=Q�'�ʱν*X)��A����\�*�O<��漃�`���c�B%�F??��I(뗅4QM��,���x�N�&���U�|b#K,q?s9Je���uM��D���b�p!���I��7\���-�ݞ�ўw�|:?��N8�G�W�)H<�R��Ձ�#^,�&���:
q�`��'!�LyC��^���F��UI���p�ƻ���R�jV�eD=��޻���B�ֱ /˰rH�F.�q�o}ɿqV��X<K"�Jzh|�>�1�� ���/���tL�l@�Fo��T[S�U���"!���M�
;S�3\�3v;80�}��K��� �����#i3,�1HV��Q@x�Ѫ��X���~�q�L���Eb� �\^0� �{$o<���R���ՠQ.h����4�4�Q��6"E�d���j���A�����G��1�>4z��:ᣞp ��l�%z�Z
r4|��=�W�*Z�S;��d9��=��d�ח��н�4�W(l�檧�P`���l�߿l�N�	(�@s���@�I��qY����������,[Z��&(MR��ձB�g����M4����*6+�Qy�ـ�b)C^��K�|r�]E�Ɩ�dd���1'͍�bT�+�r� ��"����<SD�R���O�"Ȥ�dG����©�F#����-�g��ۊ�_Z_@H��>r|��%8G�]o�RwO�/}��|�^�1
j*S[Yi9��k�A٘Rk�Q��睻�Fw����M�Q�*&��Q���Z���v�E�i@س0���F���6������ ��uݍ���"+$�[�7�(��"`��4:n��k�2j��g'�a��ҍˏO���=�8N���~������|W�4+�:��1��(�N��E�ǿ���bX������\�s�v?8:`�<�/ T�o:�_,=�Z�����'��yy�F,�fl���b؏$�5;��^��[Z�:�R_;���n`�).��e7
հi#6�'QLRO5̃��ۯ���lp
��;E\]]b,�Q��5���Uz_��x�
�t�Gܑ$b|.�U��6�S�@)ډ%u�����匚�Ej^0�O�ŕ�bȟ����K�_�F�L�� `������Nݸ�((W�A�����׆%'!{/�u��|�r`?�g5��:�͵s��@f�,G���Z�k�]+n�F+���성�����7ՎO���o�f��l���_�"\���a�$,V�O�<n���c[�>��A�N�\�6���$j��_㾚�V�B?E�� F�>HP��,����FrdBkpǇ�@��\�ML)��D��7�e����5� X�Ρ�J,�9	H�gd�߯
����b�/��S	������h����
M�ײao��!��I�'���84��SW�_�����q�M� S�6ſ�dÉ"*��k4����¢�o"պ4mN�ϸ��N��w�g��g�?��N�e��WϹ��vW� �ue���B@�����=P�h}�m郍�S���C��+��ȅ��#���h^1��j�OS�8,&�82���Uz��SfN�ݡFک��Vk�x6C��<�lmx��D�/�I�!�ZW$י��y��$0)W�$E�O��9���u�Lo�B̝�R�ͱ�k.�f;���J��2�c��#+�-����wQ�&ä��MyE��C�7�=�����Ѭ7�x��wpg��nPֿ6��ϫkL��7M�॔\L�5��m���f�7V�.��ϑ/��Y.8@=3�߂����S��-S����sLE�l# ��p�~o΢�X�92���-�X���u���yܝDU�2[�������}	 o�Gl��B!#9�Ũ�uu1���Y�Q��A��ږ���{>q�WQ`R#o�a�)~��o~�Cc&��`��`����Z��홂J�/�y�U����0�G�׏��R����ʯ�(����	��o^�l�F�x���8R���~�`D%�ʓ& DJT_>Tm�]@�"K��E���L+�[<r%!�v��9�&ڟ��W'�g(�@�xS�i�uR)���'P�o$�䕑�q`��ЮBߪ}�
,m�Q 5��H�h�����rЦp��#Y�;*�Du�!�Tl==�UC<��3䮠t:G��L�^x���b�t�E?���7�ѹ���&f�&j�$�ؒ�(�H^��M�>��E�d�B���-�-�!.�q`������h��Y�[q����:�49&���ù����� $����?0�����!�a���Ȏd�I�ӥ���Cu>����92s^�õ�HND� ���	�҇G5z��<��V!0��D�U�5��;�j��q���������T���BE��S�_3�k���:���?���["/�-:�ǉ�5����K�A`X��}����L����}�%�q���fy��2�����<�7ń&s�'�YL��o���d>j�Rm����N��"
 8X&
E�����$�Q�a|Z㝆����pZ�%���������#���~��+�/t���w�d�%��S��aEt!k}��sh�q�e�Q�u� ��`閇����EkƜl�e�V�[pQa* Y��4�����6���5��,������GY�¹l� �nS%���_�
�uo8�����8ٟ|��=�	�m��g��q6��Y�~�@�D	���h�%�L@���i�1vp����O�Kx�-�]�zd!~2��JZ���1�w�Ճ��[�t�w{��������pB�}9(�i�/��ƍ��7nHbX���Tx�O;�W��Hh��{DM�
����^�-�4���[YT��}r��'j]@9�xV���M����L����1�K�����1^����@.v��V�VZeȄkdΧؚl�Z���7���B�Y2�Ҫ8OV�\�$�
��2E`w^A��qJDz����x��w�NI�:��;�G`l��(�L-�!�%�IC ̀�@�כ�i?��Y'x�C<���.�^�\���U8K�&06ǱDˢc$��|��qB\����v����!k><O���	ܡK�d���J�9��3�b�d�c�,B���2�L�fЍٙD���|e�h+$$��x7�^�!��L��6{ƾG�<fY�tU}o��'7R
��/�ިC����~1�";%w����T������6�CQ;L�?bq�Y�1�����Q�=�e`D.�Y��Ĕ�.�!��3��'�W	P.�n~υ��[�� P�VOdm�'AP�:��#�P!NF�y�8�CJ?��ܥ�7�"H�*%i�eƏT��P>�A����A3X�V��'��	�JD
ðRF���gG-;�2|����]�'���7�zw�/��oE��>��D �M�Me�%Ǘ�ښ���v�G��_����d=EZ����ǉ�]����40	���x�r�;$8��|G�*|(�+�"&�E ^#�<�_V�?� ��?�@"ٶ��ҭ7�(���U�*1�.�fkIiؙ���{��,��s���!�����H�����g4�T�Q�����a� Z��X��$R	�be\ԑ�L��|�Z�#�,TX\m�wiP��-r6�v*�^�p��(���z��[�0�F�=���cu�z�ی�I�i��F��0��d�j5��6O��_�O$�sF-�7�G�{r�R��,綔I�T���@��\�iA��F�<�w�V�����Y*Е��޽�Ues��r��^���#�"�u��G�7��Hh�
5^O"��Ip�j�Bmَ?W�9����R%���Q�_$��a�ly_ڷq
�#�^M�i�\�b&���+��A+�w��0�t���أ���~��~�d (~n�r*aG��}l׼~u�Co#kpڨ~1XV�WJb��O]�<_/���v��㣹_`P�t���5?�
��@@�%�m ��p�c ���3y�`��à�R�y���O�^T~��+�t����=�� +�`q�)��7j���)��ڥ����-�$���xA(hOZ7*=6[ ���f�k[��s�F70���7
p�T������ZH���l���"���"c����iXh Y`S�D��Ү\���� ���q'i���Ku��R�B��4�-�Jkr�;�)���� \��y�sZa��$���qO.�zi�z)�5�nD�'iO����Pl�m�9l��\~y�{��km�e}FK�Zi�Ni͢*�`^�Ŷ(���B(�<�?W"��-'�u����V�},��5�m���	��R�ERa����{����HGq��j=�15 �7H6:Є�9J���Ԙ0�>���C�sh(c�ld�-��{��J�zS�s$�*���� W�*'_ �Lh�ށ�ƨV̰6�7|> �C@�}�j@78gD_�h	�����G9R�I@�g��'p��U��J������;�	R�q�!�%�rRAJ����vS��r�ļ�+��Б�B��D�N�Abx>n�'5�Zݠ$
�fc^�CE�%)a8���V|�[�Ը�q�.���*d>klJ�Š��y��Ka�r��@=�p���=�S� f���4!���ܛS�J�.bzA_h��G�-�8����d��
��du�3R8l�~�	�
�.��r� n6r$-��z�j��PJ�Eʰ���n���'�D������T��/K̞���
ݖ��Dƈ$/.� ���S}\a�y�)k��:��g#�oY�F<�l�� 􉁠�X�zЋ��G\���@(?r8�L�`�a,��QR�^�ՊA=��x�|
����Q�z�|�
���S±`�,/3�$���-�����:D�009��7�=f��dOY�+���y�"�Ŷ���x(#���"�ձ��j"�r���'�l�GN��=��h�u��e>A)�3�v�Ks���M	t B�v�
�LL����DEl�5��x�<�`*НR�`�Zs*�XUh��_�]S5��1�[R�(1Qj®�󔮍@�(��/�n5p��3���*8�I���=.��5DYx6���d���[as��E����n`���8�g�Qz2zG�f����6����#��`��^{]3`+�����IE�$>lη7�[p$_���aq�q�;J�L���[C�1�y�@����k�
]�]u��V�$���8��W�r��iA����k@nl4r��}T8BH��l����{?��{�(�u�w�P&����l*ɞ_��S�ɭ~�����@�N_����P��wڜ�o*��;�N'�]��f&D�y�#��g7#������xf��Z0�����{>9��6CĲ���8���]M�x���ZG�_>�wEuJ	���0iԊ3��D�΁�:�����R��=�8jJ[9�̉�M�p��`#�1��fd
(v�R
4mE�x&�����e^�\|��n6�K����d_j�"G:V�2w�(��o�G� ��Icб������zal���������W]�u��h�	�A���@��U���Qs6���C�K��M� DP.e�)x9DЋG@����-�΄��^ƾ�~��	v;�t.�uն*�.���d�ê���m��K2͝��WT;�T<1ďil�F8ý���C0V��⁈�w����!�z�̫�(%�|H�_����Z��$�� �c�"���o��O|nL�3Or��v_�N����#�JqV�'`=_gBF !����hH
�CF���c���h�<�+`35A��ƈ��c��4������6�8�Dn�O�RG��m\��3���eol|�;%2�8L|�~�ŭ%���D�Q������-"�y�V.�s��>���!`��C��y��ڬ�O,��Ρ�Vd���p�����.RΞ�(���#�-�lH�Նq{[�Q��'j�X�����.%`N�0��2�;9����
)�ԑD��;����H��b�d �[���.����X��G�v=�w���,�M�I6��*��mH��c�@!�--د�+d�y�il� |PK��Sg�
j(�{LV�+����v��P+��x��#q��}�O��N�h�2��w���;民����?�T�Ǔ��L�'e�7��YT���ܳ�U2�W,�>)iW�\y4�t��$�P��	�<�G�I����|V�v�eﹿ�`]s�ld�*��������t�ᒪ^����"]szӭ]3�;2�NkIj�)�SN�k�f���ā&�J�v�M��wk��е��K��A�y�Xy斓+��Z%�]l92x�l9꠵�@i�ݪ��V4�Ίj�<]uE�t7�G�t����8
�_L�ʲ��5�4	��MЄK"�A �����+�_�M׾{�t�jK�=�ҍzq��[�]f�y)�+�
��_�v���mlO=��e�>��)��o���T���oEM>U98�;DJ|���`n�W�7y#�Oz+n���-��;��GJ�k]�u��V'�`e��;W]r��kh�WT�Eio�Ukj: e�Yr+���� �2D�}����-�x�v����
x��B<^#���;Cs��Β* �	�	]7��ĩ�?�����ӓ'�g̅�>��;#x�JUBQa�ز>��f�mX��y�,>cx-S<̍3~�h���;�;�Fg�� p�()������S�N=��s�Y�q��IV%*�yt�����c�v�<�:��j�/��JMz�x�G�nX�����9�Z~����(`���A�#-�g}]�|�Ȇ��&J����F.-S���̘%bԾ@|y9�+� +$g�}�.�o�V�}������%�&S���vkB�I�V�Y�8�f�8�H"r[��c��#̫o	�9�:g���@D{�].@�x �ƙTYj���Z�e&�Y������Κ3p߽��|N�H9S-8e��4ʜ�L�~ߪF\��-�f�܉jx�_��?�n@��t;`��U$Я%$�;v/Io��{��A�3���5�!SXn��Z�&�.�F�e�<7B�'���Gm"�Yq!V{@�M,e�W`�wL7Y��XY�:�/68�'C���#pU<g>0�.C_N����?�DA��*��]m�U���x��d$C����jw��'(�~Mp���	-�w��O9n���$(�KW�w,9�"`��mԆ��g�����Hb�g:�@c�n�/R�T�ݪF��<��&Qyo��ܚ0:������H�󚴘cC�Wg0��Y��-��ԛ�s�XϙCߕj�I(;ʊ��!�=^�9���nc��5!�uS-�hr��Vh]�>j4�x3��<aˊϊ�u�CI�8�3E�K(�����b� ���AΫ�z;���O�������g���h���8��cK�T�A�6W�5�X���Y
&d�*���Bn��d�\p��e����!��Jݚ%�6J��Q#2��S��?����:�H
����!]x��1^.-�Jɀ����o>��k��\t�����,�ɴ���nQ!���3|<�=y�Ϯ0�7Z��Z���Wl�<�M�J�%�P�UEg��Qx@�O�P�i����bYj�ƩX��H
�J��L+A��|��jK�b|,�ӽ�>�B�iC����|B�_P#��^��v�>�ĎP���!`���K�(9L��(�����7#Ƕl�m󟐸:�O��8*rZ����BBP�ȿ��`{`<���x��ﺘ�"C�/�C�����$�H�P~ 
G�s��K�0O��Z3�b�a�Nd׫�dy����b��ju�fo��)�r��n'��XY�0��u�~VO�4R�DjLo9�N��������4V��m��PKп���4�P�9�X�,�3��y$Z��<:�G;��j��F���2�-��G�_���)�)PHG�e'���W�/�lQO��;˗�7i�0c�gcj�&�{=J/����Uߜ�{��y�3����=����J�ؑ�6:a���ď�`�
M�P�A@e	��1J�C�j�V����
�N�nҢꇦ��(	!�N���( �������.�,��,�b#�e���D�xRÕs�]D���Jo�Ra.��	L\��e?&zx|Gu�C�J�87��]�:�d=��/��~a�.#
.�(p��`!��J<����s�0c��	��#�;��M#z�Nׅ�����\��<�a���f���=�S��X�g|q���n�,��f�6dPKY?~9�ڀ�%м�~DQ��Gd5��dmM�����R�"��]T�P���%�8��9g(���b}Z�c��r��kZ��]�G;���5�_W��Y��#��Sv��q>ʔ�`s�Ķ'�����A��(�8���r"X�f���t�+6TT���y�UN���+�7`���~t��,�W�9c��,�����F�.I�ܫ�o��H���cE��/�oÐ���*��HKr����s���wp��E�i\>���@��K5�$(|�� f,�6�,�-�"��8���&��h"���n�?�kҜϬ� 쒆z�Y�C��|8�VA��[̂�7J��+ʄH0/>9�S��u;d)y; 8�wi{:M�[�/w{V��,p�\۾�N�P�i�}GJ�Ȫ�~�K��#r�ǆ�tـ�T�ʟ��챻2��cB�"8`U�8B��U��ui�W���t�R�gx�b��0�'�K��62S2Kz�!��\
�G��
#1��v��-�8�8U���<�\|>������`P�_�t� ��������x�a����U�pW(Z�?o��V�f;���bȯXlzl�Жq�� ��W��DuQ�lU�NyIu}�P6������~+{��E8�����I�M���I�:��1ˁf�g��v���C�ٌT�RXb���6�-���މ��������n��O�s�($��
h��p�E��ɂ�lF�<|����Ù�2f��[젃�"W�~�_5�Т��b�^��<�����8�b��ߚ�w\/z�P�f��^��ItkC�}@�<��kP�cST'���K@ rȊ����_�^M�Va0�^���0�*<��/��!�S��'2���W7uR�N�/�LC�V߀�V�ry��\�:4�`�RM��j̙8Qǖ�Ȱ�^g��	��gP�nX��� 8b�ԟ���5d��C��c��ն{m�+V�X%U�7b�:<��S�Cc^�p�⭸���56<Cl�鿱J�m�q���"�0m�3�l?}�>QG�l*�8xd򕬂x�O�d���c���o���R�P��?�R��������A��[��GG<� :���t�+B����KvϰqnM���*Nޔ�\���f�\Sm>��nȭ�KQ.�Ods�;�+��z�2������s��)�pg5X��7��A0��:��h�G����	��7�m����)�Ȟ��T���Y��]G�o�ڧ] ��g�C�؄�P�Rw��T7�"�h.��
2�p+�/$�$_�fٟ�<�Ck!��7x�9iٮ�%��W>4�A���ץ����m(E*�JE��Hކ�U�z��-cj��жgm�nad�qW��Ӵ��{��M��/������b߫�}�-�x�M����د���^�k����K(
��"}5����)�=���&�!3��7�J[vơ��Jg�K��<�6i�B&�;��(�{����Hе1qs�B�,~�T��w�W:�b43���'��1��%+��Jl�!���@��ˤ@�L�g�P�[����0j�Jq��}["L��&^2N#��w#�(�q�\|�T<��R�<V�|�4?�";��دT�M���#˶Rk��u� �����?��S��ҙz?J:�(�49�Xd�K���wjS��(��19����-� 
ه;L�1Z�t3���Ҿ��zҺ�'��]5�<�4鋌��𐬍Vh*�������i%F\x>��bL�� ��&�=�I��Cr�C<��d�������8�~x����M�E,��@��4 �?��������T�=F���	f����=�"�u��$#�%���#C����ߠ�G�~�ރ>�+�(NΛP�+7���~U?����.?�m^��x:�w���%O}���8�ce�t��ӿ�lF�>U���� B"/��E ��cn�B��3�$��~��}�y�A�>=�d"d��|���V����N��� f��
��nK�ќ��F��P3�i`����O4�W��{!
ɢ�=�T�Ii8w�v�������s�0�I�Ld�V�?���H�h�>)X�_�휦�93�DH�.g�֣�ʝZ�� ���"WǠ���ss!7�L��qv��Ϫצ'��ft�j=|#W�c7���E-͵U��pM/3� P.�0\K�B�݇�j�v�S��|��i@~�u$|.�Z�:�\2��[�����F���L�3��	F�I8`�K��Z6��pe�*,D��(��F�MB���;�H׸�*0{��L@�i~�U�E�6�L�~��'��?��jA��� c\$jɜx@��[΢��d�i���5z��ϐ�ϼi���p_K������N�A��ߺn�gR�����[�Z�;W��ޠ��6|ڈ�u+
{%�)�OHn���!.�b��`�JR��b�1t��{�ǫ$p����_Z��*�S>s��ߨM�d.��#>�����'3�S��}�=A��!��	euZ��$�f���9��У_l,���cJ�"�,�
���&�ץ<�x9i_��9Gq�?��#*�9��7��7!_�ƛp��)C�����9L�W��3���p���?tPdyV�<��}>/��p���Q���5�ӝ���D���m �5���E�&S�g4�2%�[2�v��?,�����B	Âʛ�,�`�+���]:NɖF�9���y^,"O~;�� .������v �6����?��?*���\3~�k��م��O4ԉQ0
�=������)p�5��lǌ��B��� q&�X��6~F�!/-=�H�w���DIyZ�2_z+�<Zz�oD �)�_�Q��Wp�ئ=p��|}ѣ:C��/
�R���D������њ�$�{�<���l��������l&#繕GO�k�o����g�1��(rKSA�ϻ�������J�yf��y��C:5`eqUp��iP�j	j�M���I���ޱ�ЁY�l���Z��̓�5�y|㝿����LO�o*}i�\-Z!����$���z�BbtJ�]1��!1pP���Ne��09<Z@�4"�O։��T�ڽ�o��!�}��@�>J}�+c8��!��'��ڸ��2C~���Y�����T�ǭ�+`�\bW�c��Z��-�C������*y���"��>oB|Fϻġ�m�q�P���|�_�/��bӏ�{X�/�O�ۧ��] ���f��,�����̓2��[	r�
r��Ӷo�����e��5)��M���O����A��:[iד岹3��a��1?sz�0�"G.�#-9��h�A��Ď;r�1۷,��3q�Ř��R4{����Y�ӌ���}[�����qV�~X���8V�H寅to4U��@�H:���·�n���O��������@x�5�=)����[�<��U�I���W�$ !�ˉP|�4��s
Ӟ�?[��轐jN��%�J��J��b�Z`��?VIϳ� ���H2vQ������[���px���!:/c5��el���A��ʈ�������~RnJS����4��&$=&�H8���jO_�rM��L�"��e� �noV�=�@�F���V{�&�,d���t��J#Q٬���55 ��A�Z���Yɸ�pC'���aW~n�KuÉ~���%�˃�n�^Q/��ܻ�D+�Xz�a��~���,O�Q��~�lڐ6A���$�t�XV:x�I����s�^k�g-OhJ7��AP4S���,��)����(�����NA���"	BHD<v>���Í�n��	�i�ᑬH�I�Y���l$L �e��./�1\kXS��������%�#n~*�h�ⱈ5�>Zr�H
jYH�%�k=:�Zr�]jJ��z�WK*�¬[����r��p#e<����գ�Ax��^tڒ� MA*2��z�Ǽ��(�3In�K_�Q�/I*<VVg;�֔�����a�%'���^S��v���(b�2}B� �\i��0^����ނK0`S��]h��-��uP��:��_�#��(������X�R�;W§�����f�5��̋)S��`v���ޤ*�{����.?��ʚ婏�]P�w�������Cei�v�ad~�6�G��Nw��괳W�/J� A3M���HuT��Ai�>�v�������"�3���`R�ګ+�������&<y@����a��D��bGr���.��pU~"cMΛ�(]��~uLa�n��^%'!�,A���C�Ec���_乡YʌȠޒ��Π�T��-VV4R���Tw^@������ڡ�#.�#N�;�n+��w�L���WG<餃,��I�~B��Z%K3��)q�K mi�I� �X�����S��1���ioB��Y>�����4%��������~��o4�Q�"LQ���bK�2���fwQ$%��p�v5���N�S�T|�0�����T��Ι���Yq�����Q�ѹ5����3"i�>�����A'ŭ�������(yC{�����E��KA��_�A�F=���T�E�ؖ\h*{\�s����6��]�	�|s`IZ]FWc���{N����^�č
�);%E����ޚ�#d����%�Ӫ/�dh'֫!���HZMob�Wl��``��čڽ�=X�����GI@|y�영Q�ҧ�y������U���8���+d���SQ�s��`꫒�����ܩ.mH� �/��ī��`'*h�:K�5Q}Cr�=2o��gF�>�-��Y�e��4�O9�~��p�}qeG:�:�&��α�G%�����I��'[�_t]A�����:�e#���n7W<ۛ&]H�lM�vz�tl�>b�m"g��/(�$���Q&�M���W^�	7�e�w�b�?��-�A�ML���K|�F��W�`�P
p%�~ȴ�3���g ��y�E �F��KNZ���n�X�6��b)m���MI.��X)��n��٨B�E?������ƀ	�	:0��q��2��r��[d��U�边����h�;fJ���?u%ʌx&��ity��G��T܍�Q��A��gd3x�m}3�'cWa)AuQp�^d�ha���p��ٖ#t����h Xn�\lbr�5aϴ�l�����e��*���al�.��`5K�RsU���(���<Fe����eXnY�����0��fV$�(�/��R>�c�_�%/��-�SQ�y��.�폟��'NLC5w?�)�#���|�4�g�>$��4u�����W=B���H\f��K��.g�)�>�5�V�rK��Q�8>��#J!�Z�:J�m����̎#n��\:����\Q�ӥ��h I�CN������R[��m�S��)gO7?���	o��f�xT�N�Ķ�I�qKc��\Қ���}r�q.n���B��Ҡ�?�&�Z�"��ھ������U�~���.ݿ��ՖiOf�2�N>2(U�{����I�^����#&R�akHr�Si�=\��tJ:���rf��R����j��%�*3]<j��<"�'�j�}
Īv_��")��i|ǫB�|R�R����S58�C�#�	Rn���`S�������0�»��L�(��I[�(ϴ5�H�m�U��5�=Wf��y�ÅPyϿ��s~p�<��g:t�VQVF�T��-��]N��oy�ayƚ�H?��MZm�gPO����� �]�k�J�'���m�l֬�j�_uG^�fc46̑�r���ل5���wK&0)X����A���1� �6���1�p2�V��CbGk$��$}Ьk�cq"I��߅�M��Z>[�?r�b'{�3�.���l}Mrfds�����ߏ�4z���"�x��ɫ�~�Q����VP�>b���b#��/U/~j��D+���[��8D�#����V�a7��-D����1����|��x�f�O��ņk�]��צ;&�nJ��.F�d���X���H�e�<P��~�\Z^�q6lZ�I���<G1���Y�r 6��v�����3���5}�����5�O{o���HP�K��1��M��҃����E�!A�{!^�|��9�k7��W�:�N�M�B�Z�L��*e5=�쫯�el ��dI�/��FD�r��C��*둥2B֪�➨G�|y�<�L�Өq�b�t;�F�j�͐����K�Y��'��Ar������%��=|j�d��5G�Y��H�m�7��><9���6�!Oa"�&^�r�	9�X>����V����~���\��јg"�D����[\�9��S��;��Z4 �!�A������`�>2phE�d�+4�s�>k1����L��$ip����͂�5T����}�U��5ׁ��U�P4���Ꮁ�ک�rH��WW��{a�*���e\��9H�����%&������^;N�t��V�����#w�\�B��U�61ҩ�-;'�A?.E�^"-iNӨ}s�K�K8-��"��>:w��-�b���8�]����G�-Q�E*�9�qv��Ɂ��+�����3�2G˷�7m\��Y"��K�T��Q}0���l11_,K�Ȓv���)��o���!�/�c$~ҋ��#�r��������9ٝ�'	ݽn�V�9��7�o�4F��Z�`Vݐ�B���7?�#غ\�4�ʥ�����F�*��rw�J��KdWK�����x�Pj^��J�����ĭ���έ1P)h2���d�j���n�ʹ���O��� 	�pP�m����>G��/�C��A�Y�W2;��� ��j�K;~m���u@ʜʲ�t���ɡ��R��̻��ϦN>�MC�2���勜2o���m���1�ݶ#+�
�K�|�Uǵq%uv�gJZ���ۃ۸t�����}����#���W�!H�WCy��?V3K[M5���Q��N�`�i����dB2��!Q��+`��;d&��B�����L
?��*DX}� XgVҚ�n�0z���Nw�w���K,|e���Y���)�|\��_t�3p�q�Q|/OF��7]��Sˁ��TB��������t��D���8M?��]��,�]:eh�e����	��V�d@�>:�E0]��%4j���Ъ�b�3���9Yס�#$&��63�?���ݳ��7�� l��簢��]e�@B+WB�� ��nq�)��C�dn��!'�La�C�	�K�bO�������C�5� ��<�Z}�1��W}�1��I��Mϐ�@���5��T��Y@���^�_~�l��r�K�c�~3@sE s�$��HY�JZ����<�6�+��
�ד"��6�
�1Fa$'��-.���$��yҝ�9|d.�_&Qa�b�$r���/��%<H(}��Y}��6F
�I` O_=�����@�� q����gs��~��3h ��^�Q����5�
�l���yH�]6�Y�W��}�&��?���}�-q4\�C[)����^�V��ܹD�3�
]�uR�,#/ڃ����RH��.LY6�D����>��Q�����e*+���`��U�P�)�r���@�s�Igs�5UV���[�o��{'ڶz��Fz�\89��5j���ce�����߱���i���21M5<�E�t��*�I�k�K�����n�l���e�_��܅}Ǔ/�l���ܐ��[�!��X�{05`́��oy(Htyk��0	m�}��^�*��.[KEAx7�=�w�r��~x%]v/�}�?Sx��g8/(�����#��UH�%�Q�d/2{��4z=Udr�Y�����x�r����Ŏ����ߙk��m��π ����_��J��ޅ�m�r���sG��4� k�r�A�O��*�@fZ���)�=����. m�<��(��N4��%�L���� ���x?6u�6�m���:����5��ɺ��y�J��|��%���;��떍�RG����b2{>8�-�m0�I.m��(�Q.l�
v�T�,�]��fK$�\?�uj�X*��ř�O̂�W��Q�����?��V�&s���Y��QO�84m�����V���Mb&{,7�'��TH�y:������4��_y�__/x�nV����}�Y�FQj����,'vBxK��M��R������!��!���sZ�ۿ���_�jpv�I Y����6\��a��3��]sD��F^ye,�Y�%.LY4�  �A�����W������v��Q���s�:B�nuS��b�ܪD����,��u{
�S�o5j�x�H6�	q~4�ƹ��I|E.Ei��.���'���6��B(�U3$�Ɇ�/���#�d���~�Q�XC�і���9��,����� 4���<�n���K����� M��dq��!�v� Y0�hj��K.������*�¤0��ܾ�SߣѴ��$Iԅ�d�L)6�U-�n��1�[�T �ˢ�^<Yy��N9�Ż0��A�5-���V�Q�U�^Ɩ�b�N��rVr/S�Z��5�͎h/��g�oKX��_�A�����3Uud�L���`�4��8ǝ	䗠 ���E��M�s���LJHzRn��_���4Ҽz UHdX�p
V^ln���q1�;��R�Xx���딛���J̩nÎ�\�A��!Q_<�^P��[���Td�Q|��j�jx��os8�H0e�R��k^��>$e8"V��t���`�����֝W�=���\�Z'`)��{����«F*P(z��8|�@1���YI��M擢����wř)F��^Y��s�oW�~l�:�eq<n��$��C�^R�_���p��%+�M�h"��B,�cb�Y�y�_J@����#l{�%�y�l�\έ�๶d5�ߥ��Y��i��׳XM����|\�j@�d��ü��cn��7�@ԟ#����I~��߰��������V>���m����s���"�+�U��@�
�%le������:�L�bFjs���
q�+qA����+�!n7j�úC��j�mn��b�v��D����L���Xw1�v5A�|�Ĕ���b`�H4)�K&6ÑI���S>�؀�� 㘭v��\/`�$FU�V,<�JF1�e�7B#�ثH?��s�����:	�����g��P0fu�P��]2�ur����^�F��k��$^~��)MC9g����Dή��"�C��j'JJ=i�Bw�{�㿶��Ny ����V,���m�eڒ��)�["�걉�,*P����Q.v�o�~�L��4����� ��`�ɃZ��#���*����Юh��WRNǮj��7e�
U�Hq8�|���qǧ���!ڧj��\�r�{D�v���L��{�L�i�E��0�X��ug�|{&]����[������I���g%���g�Gi;f���[�P4q.eH�׋�Ѕ��|(2b�����+��h^3� ���zE�e� ���dHM=������\ْ�5�ђ_;L 9�|�8�2�±Io2�mP ԗ��5-\�J~];����E%RH!�A"�e����nq���j�a��r\8MD�<�ô�@�L� >��A$=�� OӔr2v}��tM�Ly���N#b�u�K`�}����]MϞ�3)1�i��H�^V��T47+G�xV�{�N�uc�����"N;���_�)�8��I����e���Xk}��X�т�-��I�f\!��"�i�%������W�Y�1A�����%_��x$Ѭ���f��|�-����u���7�iD�8����D	x�|�D�R�s�T�m���/?1�~EC����DTr���O��o�U(�
c�i��,���x��.��(4(ۦ���{2���Xr��}�P������K���M��(Bϖ&����E�!�d����!Ϙ��"��o�D��|��C�ͮ�ֿ�AbJ����GY���������/)��вk��&2D;��,IRQ����B(sK ~���>����!ٍ!�pcf�7���ª�	(��j�AA��[�����h�̺Y���&@PVŘ�[`�80|&��Z��9�]D[�u�-.u�W�*�\n"�B�@�����(��ڲ�y3&Hhf����f>|�7�Mdԇ~B  3
.�,�}A��*y�Հr 9���� �4T^���9�%e�"�a���b��zW[���r����!���R2���m����^��\H�3w��c+��+|	�T߬�Q�Θ>d�e<ઙ��6�*�9F����	y09�o��@�9)NxƦ4��K|9����5&R�3L� �a��]�"]%�d`�@�S��x�ӷ�n/pY�	[��>�]LZh���WF2��(��j뜮S)q�s:����%q�!�U�8	i_;�\�o�|
����3ݎb��%���p��s�k�t���UOd'l	P�i��hȴ a��Y>�ylXud����gn��2��u��ňT1+�)b'�K�|�w}
��f��M�7��\.z�z�p�;u�w���R�@lW�pIK�������`���/t��Ԇ���,"5�H���	�4���=O��$͢Bw�iw��m�noeެ<8���vê��}��!M����5����B�T��dX�~�u
/�G�.}�T0\�.O	^]��(��_8Wc�ël�K�V(je=�Aʱ<�0m��$L\GTt�[�_���<C��?X���) '����'����.~�u�1+,��ۻ\�b�<QHAݮ��M?$K��X�:˃ �=8i·�㐠~!�lX� �	^��G���"\����HR��aM�&חA[��)�	�[�1��^��pL�%Z0�Q �Oh�<���R�k�m�֥�A�`�%jxH'(��;�R.��=YV��&����5�;�mT�Y���wX/M�ߩa���Z���%8-/?<_��rлO����(�hϙ�)�0���߅�,}v�V��a�n7�y�������i��l��}���C�l��(�$�_�c���}���=���e�|L���d�F�rӉiy��6�C+���7U�0���hw̌��X��vM�b�]彲E��?i�Hׇ�S/|r��;��0Չo-F��[[��B��ӝ���&�k�/�-��"pI��.s6#�x_�pi�yH���J�~�C�f�ꏘC|�b 		QGmn&Z5T(���,N��~� *wɝJq8_�U��k�q˳��Fo$ڂ���6aYT1��L��,Q���3\��6���h�W�D�a���mG��	e�(s�9aв�5x�����e۽��xL�L��`W-�Bt���n�������!��95��e��̕���zc��a0~ �T���-�Oc�����[;�z;�-�Y{�iK�����+}C�mޞov��\���6�1����O����[��Do�)�^��M��(��8?��8�=��_;O��y>�3��E��Hh^a��ץ��٫�"�S F�y�]��ʳX��Y&�Cp*}>uZ˄?��(g�ZS�jVG��I|�'ED/�i�8�f�&��,J�&��U�~uly�ƭ"t�*��a�GBr�m��ׇ,3�%���[S3�b=�V%V�Q�jќj""J�̈(�Ā"�dJxUA�$�3�����żC��C�J36�z~:�V���QI���T�j�w�/mn�.�^��]����]-�V�{�gb��֒��34�� �0VӷJ�ͳBVʜ@[��I1V��\,�B�v^�|�w��e��Uު�D߿�k�Q����|�/,"�����&�+�Lg�@�dw�3������r�z�����.�����T-{;믇җ ���Ս=���knϸ�b+��� ���)��];���gW�b�Az��v% f���$��쿁�MI9���'�.�/z9 ��"0{%$�d��C�����W����u��}R!H?�L4����?֚yΠ} P
�N����j�t�5E}4���qm\����r��σ��TuZ�MY�`)�S{[̕^)0t��@��&����n��`L���_�DY���{ٷ;�!��鑜���5l�.��!��_�>�kMR�)��R#ztb҈^}J�K��~,'�8��"�R�c�#&��4S}��JA�lR��y�+�aO"�'[M �Wކ�?T�l/�(Ж�-�M\��LkP���/w�s��B����Z����bk(Yb��s��ޘݱ�=�>J�39�^8�T]�\��f��2~ċ<�l ������cg 8��};���坡!!f&�����@�tP�U8����Ä�'1��Q�Cl���:��f����I��5�4�'�uȊ���pc9�џ~��i'�3K��N3�"!l�FP|vM�h3����x�3(��AFr����6Ke�?7TB鋣7<;>��ޭ�72���_�HC�[[�z�q|'���?���O�4��l�,�&�� �/�����Ʊˀ�*�(��}|��BZi�����K*��~�t�Ѐѿ�Ss�&Vc�|�u;|�ErNY҅�����v�qL���+k���@`#��p�͉>o3������þ0��;�D�3mqC�p��=�v�
��O,�;E�b�7���x?Ȁ \n�۝�I�,/�U��O��|F%=� $���I���9}J�KZԔ�H�7�=Ⱥ�Ey|	�����aFa\��[����U�?.a�Z.}�N��]'D	x��[3R-�x.�&0>ޅ*CZɈg����Rkb��1f��z��e��r�J�G?4n�ߊ��)F���K��z[p�!^m~ȼu{��.��mk�����2�倫��Ŏ5��}��o�N�!�g��*m~�n��+��=eظ�o�'KT�*��h�E�J�o�J����+���E������0.*lv�-��Ã�3��w�KsV]�һ��@>lO�@A�jf,��nt.ؠ���%i��@<�2����B�!i��#�)�7�I�&U����!��(��P�G�-��K/u�)��IԟW^~�Յ�S�ߺ��}�ϻ�lYO(ۄ���"fW]��]`=6>�]ʂ�JCENz���C
�򴠶���?��T�<$�U�� V0���{�xx��֏Z#g+��@������R�,n�Ԧf���y�R�]��	C	�2ך�ҴH�^�(��]o]�:�#p �[���*#���iM:jĹ8��(�B,���ٝ.ғ��J�ҿ��PsNf��݈���3>�E/IoB��� F��#�oE�#��i��p����9x�*ns �=F����ENș�=��ǎ!��0�"�o����>Q/|�d���WE��(7K�j��k�t5�'�X���U,s��H �*8�JEcFJ\GW�P��@ &[��^G{&I$��.[�����=����k���q���0����S�X��C��w�$ ��1U�"3���N�3p��38
��H�����E:C�,�&ߪ��c|���~�����g�����pIY �!�{^��#��㋜b�i);0Z�C���%bֳȬ���$��
d���<��b#��K� ��$"Y>ÿ
D��:0>�;���qx������
%e�N���g�_���8P��H�\���\2���9!S\�� 6�� G����g�P���yd���N�s�U������;���	U{��[�ކ����� �	7M�x��#Fq�u��\}*>�u6Z-~�~}��U-��6�����j��_ye��V�=����x��Wѯ�胤�@BC��/%�fR�QF���$*Y���� �^r�8yT2��"4����=?�rQ�F��� ��,k�ȉ���d��O ìϦ�ŭ�@�d��`|� 3���ӝ��y�a��d�-UGQE�}��2����ޑ@BYC�=c��t6��s��9"����-�����`?
�8�Nr�J��xF7�x�����>�~)��r�� ��?�[�37��B�H�����nL5�X�0X�:GG#w06��2���=Y.���ޟL'��R����P�C�?=���
%��p�X�L�/,M܏�}+���ل
�D���A����P�~�,��j�Ñ8�<��������u6��k�E�{0t O������}�p)%k>wf���ԭ6��4z�
{k.������f�==|d$w�P-K�t�~�����Tp�Y���of���x�,H�i�}����Q	��Ip3���$Pu�&j��ن���h{���"=T���t�*R�T�(���KTL�<^��#OpA(��{ļR�jk�WA��^��ac`�k��ŉӟU״�\�N>:�0x%�	z�G��Y9�B�]��X�_�].<����!�UQT<H�_э0Yڝ�@�G"rA+�L�%�͛Kv��p&�QU1!������0�sL�K[E�^\�`���Ԝt#o�Sp��7w2�5�}� y��||�% ��<�f����)�m=A+����t�vA:O;M�k���F����u�
�Spa>tn��jQ}�a��}�DN�m�F?l#N��Y.d����Q�ow���"�0�O�U6�i	�t��&EG����軁$-��>��.�&�H>~ L�bR�,�Ļ�O�M���hV�[TT����"�ӑ�*i������9dB}a|~�q�Ns�D{P��_Q��>φ� }�/�(t0���9�vѻ��+u\F�)ns���gW�KQQ`�*7�B:ΗWu�]Тl��ǌ1t�ݤ֠M�����b�q�����99qq���NK'�Ѵ����^el���K�Jbg�s+���s#AӨ��+{:��N�TYQ�*璚#,���[��K�ʂ����n����\K�gOx��J2�n2�V�'��Äz�7��n��m4EZbv��,B����e5W ?s�̀5&|�B ]|2T#��?/<�?��m9*��{�#��Yн�H>#w����3���Tk�N}��X!`U(�?�L>�����$�6_�4]��ihk9��h?[;�U���|zj�w0H'�V��I#7�f`�*c��6�b��"nEl61�w���5H��y�6r�w�3w|h�����"/)*p�����@���kisx�1N �`���řN������牡����,��a@Ӯ��S�(��!j~�2ܟ/1p/me���de��ľ��V����V���𻱑h�B(ncπƺ0j�k+L����� ^1��c���7�E� ~�"�� R8�F.F��\gV4L>�:�:�D���~K��_���z�␵(�(��0E�|�r�%P��=g�hV�`ڊ��}/&rɺ��
ཷ��#1��$�њߡ���p�T�vN�.�G�	�Am���.��A�A�toe2t{�\+Yj?�>3�S�����ԩ3ӛ�W��T��qU
x�����1����69�d�L1d�v�/�]�NT����8H�D�]\��i�:(袘�0�-��AD�X�
!�w�7�3�#Q3ι0=�O�_�6a�pܾ�!O4��~�uR����L�
�'�"H��}|u�K�7��x9k�T�<�o#�
���K~�|܋��1��ڝ%�j.��4�`����E��wfv��E�$�!$iU��(���MF�.{��!�(M�g	 �[�)V��ʜ�D�y��_�T�_���=��FP��?�!�*{���T%�y�P6�1!�O�����ƒR:��.���۪a���^9Jh�Ql���)òǙ��1�-N���L�����(��
:P@�u0
8���H�lG���g����'��i��h^j풞��}y�xb|�z?!�U6M�;����؇���1^.�-n:�{�>i���M����_��r��p� �QP�5�ǘ�b�t�ZF?!`�A\ܨ�aCxrn�Uɣb�Ck���L���������P�������-�P��-���L��f���YJE���j4l������r)�Rgĳ�Vo�u,�؈�E��!n	�.�����_�q�G�l���;u���$�X�*J�5B������V?�Mgi��V��={^K���u������X�����Ԍ���W�h~��<Ve�&(:�I��LJ�^볡n	^.��5�a ����!�Cݾ��p���"�b����Kǲ;g5�]k_�D�!TG����m�H���YT箣&:zy��C,�!�?rD���㠋
��J{<�}�ﯾ3]�`�P-���?��o��fʽ͂���^u��Ș��d���cD�Jt��$L�z�}��c0������;Z���/ H�Ne>H�^��xS�}v2Y-)&����15 �b�&�H�[1k�@�@6&�_#w �Ϊ1�D�N�Z�ff�n��6���j��k�A�=["�5f�ŋ+�C�]�~w��Z[��G�!\O%�x �و�b$A
!��p�?w ��¥
	�m'�/��J[�j0��7�۞�$x7D�PE�N���n��m(��1�jY�H BN�٠yudkrcd(˒l��N�n�v���"�Q��!�w��mpy�dy�es�nh!.����_�E.�=u�~�(1傅��I��|Jۉ���Z�w=�n��>f�׋�������VNqs	28b��������>#�թ��4�F!��_��kي>0�HR��m+۫{�c�?I^�:�̮xAß#�L~�$�0Mл�:�/�p���jI�1"�sM���)�N��LId6�� p#���/���)/hF����&�$D�:"#QF"��]E�u�ŦDo��Lz�1`;p��eTM����y� �woH(j�90�a�)�$4����"��g������[P�V����6���W�:��47����50�N��<���-��*,I�(5����dk�w钺*���Y��]^�v46@�-xF	mnZ�M7���,g����i����k�W��?�aͰ���T3n.��u"-�N�C�=���ve�E�
|���3K�f'��c ����gN�t'b�h�k�o��M�A�KV�;J���v��9!����W1i�]C#ŋq�䬟r{[%>U?�N�j,�ة��[�p��������:�r�2�|�u�jH��M�_��@���>�&B��Aݛ�d�c\&i�"j�$,4��6��0@,���TgX���f$O(��� #�ܿ�+��3Q�-���bd���!�r�ʲx���:-Ig��3q]�W;{r�iTj���1,��B�o̜��B��������?z����q�wQy� ��i臽�B�(�(&��~��-��=/?�*�+%+��@"��i���d&F��N�I�e�J'��7�U���|�d��q��d)n(�"�X�G	�����Q���h&	��W��o��%m���r�#-��+�L\�0�l�p���o���7aa���.��e�R�3k���[7o�z�H��kx�df�=�C�wG.�U�&�ճS�H�`D��'LJ<V���<!!ˮ��L��'Wjw:��}��?�sȺ>F������,�owJ
�>jQ�a`g�<=���F.&2p9�v��{�d{�w�D˱�pܟ�Ԏ��X3?��ƾޡZ��N��%Y��z��s�fH�XS�@m�Is� �g��]�v���@�Զ�@�5�DY�>��xi�[PI�/&L��Vץ��N�&R�"ǰ�[����43M@��n9��I�o��� �nE��?m�,���.�X:�Px�g�0����`�����~��E��E��̮�#?bf�pY�nt��5�t�r����o
ȃ\���{H����2)
����@-U=��u#Ĺ�Pc���M��bH�x���Ղ�@J#��W4?�	���w��H<0g/r�E�sgL�U�uS�b�'���q����Z�i��4\a���}v��]���iϴℍDߦ�҈V�p �b�601��6����S�SxF�c1�q{0��LKO�.ZB�R�&���֐�R�O���a6N�W��on��L.aj�th�%o����/qMg�[���.7����@��/$т{tpj)���d�5�Oo˰�O\0�EmcH��t:rT��n�KIm+ί�y�:6;��z��p7�� �M�"�F|��@fy��8c$2@����{^���b�RGmS�F< ��"��5+��5��]�Gm��h��+�=����;�cA)�'L���Q'g�� �`���p��ވ~���}ds�1�`F����W�P�͗�3�pv0Э�v�
Q�쒗��&^i����A0� �P�s�0�P ��+�hО��>sz���ף�n�>]��9�ɕ-��t�|W�����t=q���2Z�
�G�g(�o�
�#%%d��Z*�K�D6��k����Kd"��O�W�ӮmQ�ZCl�1����z���J�ڔ�3��\��q�a�(��|x-�)�AKJ�+hG�١�����w8�J�փوsr���o��%cy��HE��J�-��T�õE���J��sG�fGLDӛ*ٞŢ�Ϙ�	!���ݳc'p�1b�R��J;���T�� ,�Z��>V��w�\�)�W��s�����	�I®�w�O����oX�6���(S���U�E��\�^���7{ר����d�vl��	��X�Q�B�'�<��}U7��o���č���|��)V��Ј
y^�g��l�t�@-�&e1���B��3
��W���� ~(Ls�Z����~�z�iFz��mF\s�$t�?o�<C�/9�����S��ۉC���qO�*�(I蒼?I$&���m3e?�B��U�e���v|]U92<�ř�Ӱ�v�l�	=Z���@E��k�2I��N �+6�n� K�2ُ�l߁�~�S.�S�-T�o�Bj�Z�bX�f1ک�QS�I�yy���X�lDJ���.��M���tK������Eܠ����ko)��6q��5��3pWhw����]���؈s�i�����ʍ�~�<�N�����wrd<�!DU �S�Yц��"E�N���cRd:sW��7+����d�c�"rV-�б��q?�� g�I�Ȇ���	��d�f�Og�j�mF�[�2lE��8�=ML"*��?@�:�Hx
�?��K�k^,��(R���������:�2�]�����Wg�&j�����e��_�I�G�yf���]�j��命���yaW�Y�7z����p�wVK���,S�X�t��8�m0o%ݎ�� ,���YKV|~;�a|�B�&k���F��m�����	���Ǯt�I�v���4״���@���v 58�:tS3~��[j`}��g���k��8�eS ��t��[�::�������?@8�mD!���`]�BX�D���9pV�d%��ױޑ�r��! �ћ}'@P��6�W6dh]y�%G=��������~ZV���7���pd���ﻑ:�j��h�R-Mxz)�R
,��AŒ�MeG�1����9ѿ�4�M*��I�[��MD��$#O��0(6c�L�Rҳ��R��_��h���#q0"!#�x�W���%��|�܋ei�a1;�"'�т���u�p�r5VcEk���n���_g��0Hp�ȹ�b��(��%:�Ef&"�VQG�+X%�r��ե�z=-�&�i_H����Y?yΉ�����Q�<7�Rϯ�j5����t��'�v�zĶɇ�������E��|z*{?ݖg$j���� ����hQ��zsm��k}��A8������!�y����r�a��l9��ʽ�B����Ӭ��A�Bd��.k��}j���}�*�]�}N���e���_��JE�	��t��ճ�����"m��;�T��J|X�,�/��=6��b��`� I��Z�o�OnHE�R�Ζ�@k���+���x;��5g\q��{+(�Eg_X:.��CZ#���mS]����1�e���͠�ѸD���"_(���t��{4H��N޽�?�,�nR���p�H��%��d��C��S��!��S�	�8&�d=�v���Z��N~jᗬ�W(�dQm��8��~�'�������9CAZ��~c �����2|�!)�Y+U[�CyU+FB|b�#�y���X�0�8�To\,���\e\��>O7,x6����ץZ�E��*�D8��nW�,JB6
��?�ɖ	"�L�JϢH������ޥ:qӁ��%�#b��V�Zy�z����*`�pUW��Fr��cY��ʹ#-�Z�F�wJDH�N���|>M��Aҹ��1�+�s���2A��E�'c�(��]��q6��j�,;�GI"H�Xw��M�����q�M�����i
3"��Г���3�R�����y5�u�C��6�w�����@	L�Ջctj��V�X}O`Ai� �+���w��f5�w��A4 ��(��:L��O�]�:�'�x]H����q��>L�C��I���"��Z�N�>]Ud>�a�f�mFb��7\t�R�f�6"�]D� 3	^���x[��K��B��coCi�AV���]��:�b��#���t����Iu�EV���+3R[(c��:x�2� ��H��I�#�L�MK�F�+��P8��Ș�I��)#���zo:��u��y��6o��v��8�8�^�{�C���x�����f�r�en��9MDǟ��&9����N���[��5��; \ U6M`4�������Z̤?jZ<�v/v��Y{ޤY#I�����0�tWFOHt�zu�;F$J:B��7��,t$DڗX��c
�T�X"�O��T �2_����"��r`�X5+4�SCS0f��*�Z$3��ak�f^��/-�ci��"4���f]p���'T?G����t�\J���������VG�A/6�)]��Gl{�+��U��8@�#&燃�\{#;w)%�#m6��̗ۨl��*q>�p:�!=:���Ў����Jg���j:��'q�LC���!J��#�uj %�#1��(u��pچ��6ht$a��Mh�8�-�+ �nK��T퉌��rI��i�#�@��[��~�8���t������%�h�й����&$Q�iӚ����!~L	��`^e���������uYNv��Dmi��4��Uq�4zq�s�(�[����6�o����(�bs�����ob⡌TJ�Xw�aO-n �R������&K�n~�9�W�Ba%G�pG������CZ̧s�t1� �á�w29U�������Z��5�ؐ�q��7��*�z�L��}ڔ%���E�0�r� r4�`I�4�_cܼ@i��ڣ�����<,���IO�	�R���]Z�u���	�	h�b2�����q���~��dE:�U8���G���u���������5�Hy�$�w9�����@��$�Y��|�L<�Α�Ͼ}ov��̜u<��]l��?�M��nA۾q�c�qsa����/����N�X�pL0�mE	@�ajs�1�b�����z{��CD��E�7y���N=�ɹ���uT����.�-M�M�+�i�^b���N����p
~���Bc���+/���20�9�	�T��tBT����k�O_s�"�9ٖ��Ų$%6�3�*MnU�dI�FF���������[���_!���<��2J(�/f!c����C�Y�A_N��P`>�6��h�˶�V���w���6�	��0kDٸ��́���U?d��FmY<�Dv�1&���bu�
4�f�����rt��/���mKh�~wmS���)4	Ose�C�\�=	ܝČ.q������,����� ����.*�߁��7/���{��$H9gEm�[P���̓@]=��x�jXy��$��$O[�'5I��f����B
U�7ܩ���FT�� �ΨY^&�t��m����r��)��o��:�RW�؎9�:0��i�T>O���NjH�ñޕ���h��nX+�%(dd�?�n�i��E^h�'�k\_��#���>��ӜP�T�AA�ju rbZ�V$|��߀/�H�_���M&����չ=%��)pȌ�Pd|)�Y�gP���D�m0h����0ݯA6�bMOa���8�=p�֢���-�=E+���Zw}�� sf��x�t�d�B�QUg�2%�TMth���>U@�5�~��N���.��˗��<�̡mo8�'��Fvzw9g.�Z�ǒbI8�+��o
���i��c!N4��j�jB�̴݃\�q�Q��cRK]�4�u���p�P����.�C	�EɋcLĮ�O��d`*8O�/�	/�°�^�0��-�*����/ꗄ�[f��yPU�E .F��A�n�l�HJ�i^��H,���2�aq}�!B �� "��ʘ�ѣs�9/���:��L��Bl<�_5�)�"Qǋh.[^ry�u�����)6���!F���(�����k�����^�s�T3�LO��{0u�w_G���t9�/gn]<ʒu�>�-�>�o�4�c����{̗�0�_c��U���p�-�*,�>cu���1�X�Kq��*���vY.�Q��r)BK8�D��-N��P��z�-SW��� +���uۙS'����=���f�Ks�t;Ć�7���S?�A��%���e:\$'#��Z� D��n��/�_Yk�7B�m+U��a�#��ұYK]�AWj��=�ZwPLs��Ԍ~��,}P�ñ���_��]@�Qc�%A�j�K���S}H4�����/G���C$�4D��"*tꮊ����� YIz ���+:�;ĝ�t3%���6��{]�}.9\~����ꖕ �5Z�|aMK��!�ő�	z�x�ln�:�Q��F�F�SJ�Bua���v�+��V�����F�E�h%�g7Ct�r�vU�/ �Z_aS�Z�$j�� �����W�4�m��f�tTG!���}Z�&���(a�'zr��M��S���Ú�UD��i�h�{�d��[��ڙ�_p'�k�߿�����>��~�f�K�:�d��]6]�fnD�\��j���eX���خ��z�/����>��&F��h�ZSN��4X(��}��ج�͕שP�0��߳�d�ɗ�Kң�_����[s��y���z�UYo�'V�q��%���F$pu|0�&�GS@�2]|����:>��H�o�-�Ӏ�ivTw�W�� �R<�K*��{��;)h1��Sф��z=�(�r�0����Q/���z<p�h�'V�O�1��PXtJ��l]+���ئY#�K��ꁣ�7o2F��_~I4_�ݏX��6
u��.���aiF����s�a&P\w

�9�|�b7��I[��+�<����ԵX��i�\94:�FK�毫�>�脜�d-d����֜�-ſp�Vc��Dui��]O�Ф+��G����/%b�ܭ�(�#�~�	��z2W�y���"����g=X��9��8{�t�1Nm�E�#?pP��V�3�K�^cqcҘ�f��X4L�z���p}$�^����NvX�n�s0N�r�����OlH���Dϼ�Z�R���c(�ي���LSwF���nL��o4l��.u�#\�$�0�z�������J�a�Br:����c�J�قAp��Ne�S�6��OHrzI֭�La���p��f�/��&?�r�9\�[%��Ci>ĈF�S���{,a��}nT_DI�D�R�~73�� ��H[�<�*�>1��|�;-��#��]���`nv�bq�՛��޷��7���da"eFC��EZb��0�S,���G�[2�!\��ٸ[q�e$��<��Th"6���f���;�Z`��jn��p¡���%�5�;�^8	�n����x���c姐���L�Bu[{5�Ɲ��xG��n�)n�z�T��!7����F��� �F����>zP�����@+�0���wbJ:��P�S1���J��l�gn[����������Zk�潃8�@��.=�4JӬ�zKD���΋2�m�P���Z��W+y���Mţ8H���3CB�s�l"L˦�J(mD��y��}�B	���[l>u�PY:�W�*��W�@k) �����R,��ニ,u\���61M��g}�V��6X�	�}~s���ċ�B�5Y"�؆�p���i��X����#2騄/ѧdu��>�ͻ����K�Xص��� Ca&Q��~��+����^�?�rhsY�q&%Q����˓9U ��D���ښ�K��0���8���*씇��O-�}��Q#2z�?l�7g���B7��_)n��;�g��wk���"
��Y��!���u�2{/�7���M�9����]���}��m��+���BlGZ��RV����	y��OO����{X־SY1YZ��w���O}ݿ��.��e�D1{d��eNG���qŬ��[�� ��9�E��=��4����al*�du �YȜ6��GT����]�B�a�4�K�f��ڤϐ2%�5@۳��|!�ϙ��F�O�s?� !%P����6g.\}��Y*B�!���`���d�E�e�Y���!�@|u	�+�wx���׬s�#F�.2�	c:�+�_�?}��i(8_ʡ��FJ���m����)eNaۯH�w�J�����@�j�J9T�g���u:��x��5�����)������,U�?_&���5��{�d�f�h3)�7G�o-`y�M;�i0=��lf��`�k��LPh��Y���s���Md��
�;`h��F+)���{ׄF�RR����$�?�g�}WT��HL�Q;p/�\���E٬����V�j��hf�u��dā�Hq>���q'��XW�6�����z���xg��K]G*.��C/�ǫ�XPN�[}�����/>�����Lr����5$��m�.䉒m�A��|kw�GAXK��P�m��>\U��;sIZ"�;�r��joP2�d���������2��^E9�j%d�$�o��L]�qFC�g�*y�Xâ��궅��~��Kg]͕�1_Q����A�U^Q��p�5U���d�/읁=��j7$�M7:��Ip��#�H��~�v��� �����	-$�ZlQ��F��Jp�[�*ƭ�����
�Qh�����$�e��ވ�t�.*U,� ��l�I�ϼu=YFQ�Gk�{#���$-�!wr�����X��XOA�1?�|L�X��J "��i)^ꗈ�l�d��ӷ4ҟ�'^j�I5l�E�uI���dp��2�E�U:@ �.����뺛��fx~��Y�k��0�ߠ���=n@�A��蟕����������U�Ŏ��/��#R���d�*���,�Q��K�p���IcI�r���2���m�������u��=k:����Hjޢ;}���s��
���^D8J�訹����¿%�_�?�'�@�3���t>�@�«im���g;�;���k�$ ����#�ufoTw���`-4��T���R��+��.-�vK�M0c3O8R�]z-8�r%D9�P��*֠ڢS� l�5����^���\������`���'��Y�"Db#ԑf	^,��$�MM[�m2Q������Qu���۪�0�͎�G$���?�>|L����iK���!���#�Ԫ�^(�Z�\'��a����:	zҥ��DC����]C���m�vx�NR��*�@��#?������ȯ礯��ME�w$.�]�m��?��K�m&3u޿?�V��锨���n�$u^��'�������I��;ٕ~rv��yw�B�Tk� ��<d�y�&ŰI2I8���EF��HH�=G�z������ZP�/d���R�8��S4rj�%3v*��^�bd�;��j�0�u���* 8���Lst�}F
�� 	�}KsMͣ������U���|S�O��wL���̯�Z=�L8��u��͋;i9m���6%z]�af;=��F-+�X�v���.��q�IE����J���`aW��7X�do��:��u�
Ҝqq�I�BL��4Խ՘r�����yqւ�}!̷+� �觨wI���(ɸ&�[n��L�k���y��ƌ5��8v3# /�gИ�OC�Q��[N^<��	+��\왡�_�hNu
�hY��|*Br;��~���*�Ʉ��&J�!��%7�,@v�O�juM���?�(�Z��鱘��HPt��$�o�/LC�c�}�
O��7��`�A�!x�<?�8"�_�ON�0�"��c^�J�>	�	F 
�E���#U���9��0~����+�o'���l�)��;kK{�}Aҁ�����q>�I�r1�@R٬�iC�,X��5{_�^�����)�4m6t�W����δ��)[q�cNyD/dγ�[�_40�1�S|�tr���v���ԙ�Ѫ��^;%�KU���@�)��d�����h��*�Y������C-�K�K���η|T����2&C+���CG�xU�X*�h�zR�|Æ�7�͒������8��!����i|h��$�I3izqq��C1x�psd&��x���#D��ר�6����\]�1��H����t[���`�A�@4��	���w���?�'c}	@�ȴ`4F���_k����[���qNfE�1�q�U�H�;R^��.����J��6{�;H����'��������%�S�Z ���h~�ֻ���z�r��C�M��z!��w*�,��6r�L!r�#�Bqzర��i�`�rPjdCA���nQ�P��7�5U��;�<�h�.c� @fk�
rJШ�	�xي���/f�T�+���3�]=�u��@�,_�9�VZ��Z!�6��Ѷ&t�܉�[~�6W��Ťd�p�@8h=B�*6��M3E��W�ck�:T*f4d��(k?�̟ d�r*2!�!5S��4����C7��S[�Q��Eᶥ�� �OLJK"W�c�D)�@;H�q$։�P�f�,�]�p�{ɍ���e�����ħm�?�����UA=Eأ�+%�z�O��O0�_�2�o?�:�X_$�5��T����y ��u��,�R�^\_!�84dUҗ�g��ڠU[���b��M�8n8��Ltm`T���(�2�<�򐽔������뾥�P@ޙ]FҤ�l�*?��:�(�X"�히ү7�Cÿ��x`͈֔.���"f�v(��{
�-��=R�+�G=�X*���B͘����9��oz�Q�3*�y<:�>Q��>��w+fO�
p��-5>���~�w��,��h��np
x���)��|���Xa��23�^�8�耜վ�C���p��*x硁:��|��A�G0���^�����"�la,	Sn�$½�B�T���N��h�]2F_��0֒G5c���75�i	�N�xs�~:�����0^8��ʅ�ݒ��{����E;�V5*����"d���^~Q�Gu�Ӽ�H{ �R�-�q�e��[CĻ!�T�+ M�v������#��%�_��;.����v�6���*/*�C��O\~�f2.P8�/��tO;�.];J6�a�0"�pU3��{�r9�/D����J�n�C�gۚ(Zd:���DG���FL�΁���#���?�Z�7Ėx�W�6���r	v�p_��DJr��9�aI\�ţ*��OS^%�:���EA����4�̮��k��6�_��{e~~`gbc!$B�j�������{%��%���qfq.fAn+M���f�� ������DF�p��I^;}a^�m>�Ŀ'f	���y��J�UÚh�ޫ|�����P�]r�@��.�cV�Q�PD4��>hM���^뤅�Vx���c��sl5��#m���R0o��59>��#*����u��-^wI϶Ľ[
�d�5��!�V��H^F�._��eı�o*<h�
!QT��� �Y=�4�Tc&*9���N��d�+6^����M7���	�`ΌtK*�Z	�!���f���S��[�vH*PŐ��风fmy�����Ð�=�J�|e<�� x��MO��4Ȇ=�~m��B
���M;q���8Ը�����+r�{����t;��_�Fw��"%|_ .��{��[}�r�4�N��X��a�%��}���j�˭ӡ>�`�x�F�lu�!L��W�C>�l���R��z�\�8��"�U4�"�b���ȡ:n/./`W�v\ clH7uɮ���X��HϏzt�wJ�6�ԯ}jsm�5�Մ�4����ۭ"pm���aF,�;�qB�̇��KBYN�O�	�
��#��D̖{���+��
}�eC`B�z�3T���i9c&c�V�r��&�l��,�M��U���Ⓓ�v>�z��Ї[4��4p}~��r�G�����l��^&/6�{��o���@P���1�d͉pb��Qχ*@PI�:�.��d�3'ġ�Dُ�W�!x:bD�z���(?��Zp�����2�E//S��u7-�(wR�g=jFC��#���bm+S��T�j��Β{�3l�8�co/s�,LEB����:}�����n��	��Q��a�n^Ȳ�(����gV��(O��0��4��`0��v�n���z?�����
�t��8���s����u�a�{��'_m �{�Z�.?�H���0�OR��t��
괼3��K^���n$��a�FkM0`���?�m��2��o�����᩸E¡I5�t� ��.i��-y����[N&��VK�jM��ֈ�H�����\5�nz��s�p]%���L
�0��Z�쌲��N�aʯ�Y4�]K�c�$[�$�v�&�F�`/�(��̛X�6�G+#/��g��4e��`� WHKش�O*��Y����^��A�#@�;�Qu��U5�;�*o�x�i��[	Mv^V� �r�r��Ym�~�FSK��\�uŊ��1G~*�p-�n���\"��t2��z�ۋʧ����{�S�j�T/Cj�qI�.�"2�)T���t�C]&x:
�F�[��-372�BQ/G��ʓ���Z�T�.�b�gh�v��ԝ^Y�"��G�,���uoeӦS�&xH:�U#�0s�!!!�)9�g�0k�`�8���[�W��H��ʟ��Lt�����n�3�%�_��X�^70�1%��f,����D�F9�G��
��"B.���4���mg3�E�V���#j4E/�ۍ��O�L|a��������#9ӥ�쾫2�p�}o�Rv��9/L���(��i1%Y�꾲S�Z �z��ţϨR)���&�r�CUKY�ZW&s��P9������Wb�����MG{$�@~ �p�_K��q�q�{Ϥ���& H�~��J�U^�㚺���7wɶ���)��%2�����<��iY���c���G#��K5��2���a�r�H�����R:s��Î�q\�Z!�R��Sn�`��$���O���Jc���ȅ@,����_�����Z;�l�~�gļK��r�!zg�;p�B��s:���MJ�Ю%��d<yy�q>×��X�9�zR��/��+u��3�j�1/#m�Υ�� W"�I�v�*T�%	�M�DX��?�.#̋X��ٔ������[N@T��ڷ*��#��J���5�?�l�u1��\��L)����j�F�7������K�O"1�t��|�Vac~d�T�^�ۣ��4�Z�hP���!�41#]�ЗÏ�1�b~@W��*IT���p�N2���DR2��m�����[����WZ�w�ӼN�m�UIN?W6.�6@�R����e�Y�9I�]���q6�]�����/�%z~"����r�c�BY�V��$�4O$P�U�bӤ���LN�6���/�k���qh�:���A�z3l��t�K�;	�{���S��R5Ao}��ڼ��ɔڴ�S�	�z��L�v��.}�$"� K��S`�ܷ���.K�v��y��|w���8��I�҉��b�s�0Y>0�������9bX�t�����e�ye�~�.&�2)��+��80�=����ag6�y�y��l���,e<�Xz��de̶�7�W{�����v�gp�-��He0�H�g��7}9X&�����f�]]��ૌ��c�WC�c`Y�}pq9mc6���聭��jK��V�����d��~�\	#������_�������ˌj��� �y_�yD�đ��	�1H��nf&�l�T�%��ETɩVGX����L��x�i�*���)�X����6 i��_�m;�Sl�|`��/����*�t��pҦ�<I@c�!�	�Z�N�B�k��MɱɁP��ڝaJ���`���D��l��4,7�DC5�SY㨀��D�vz�&����_ k��cN�ɴ�?Ƣ> ��Q����HR}��+�m�� (��r���ruQ
�:���O�Oxs�\P�aV��l{���������Fz�6��g+�-�� 'EY��#ݜ�@�{DBd�|�,�VŬtJ�T����_�d�U�̩��"�L��$l>�����C�����a��9+D�~���ְt_a��	����g^��ؓ8���]~�!8�E�%l�+;��]@	����U�'�W�2f�i����g�K2b��lV�#�|�b��(F�+[/����bO�;�޸�l�����.%1#�ܳ�L}��+�׌�2Zb����͍`�g��rLP�J:Q�v}���; �&��(�r�wR�m:#�
�����<K{�pC��C�6~'�[fML~G�������B�U	����`��p8G��2���1P�/5�w�>i~���P���%ܷ���� :~����u�U�v����ho�����쿔�u�
�z��	B]@v�>�-#��X��[�X��+�ERh�"���_�A����V�����<���E"}U釯V%Y4��.ԩ�G����;$�	|�Њ�]d�7��M:X��ʤA%���ޖ߲��Βv���a����Z͛S��T�kH�2!�_P命�ݧΩ��|Zr��b��I��o㚜�o����o���q<|��)M`R<##ZR��vN#�jH	�0��O�`e�Xlp���Og_Ī�޲�]����>iSS�y��,ҿ���á6� ��������bfB>T�,$��^գ6y%RjoQ��p� ��E������v��B�9[ߛ��#�~BI��|�}~j	�<�?4�Kx��<�કʐ(��@<Ca\�s��.8��Ѭ\V�\^�%5�ސu��AЃ�LU�P8}xCA f�[%��p@Ź]��K��6C�Aۅ5{�[5�[as?��ȝ&��\pȨ���0��^�5��{?`�?,$�E��X�1#�߀�eK��vo感
Rah�������h+0�z����:)Y��,����86'�����v���%Q�l��U��)�7�_^������}��\�^v�˷DLt"�Mr��	L9K.�v̀:HH�j�P�rT�����]:���NQ��L(GF��-�>�"v��x�၏(X7�U��*e'h�W�{�>8K���=�L6n%*z�`�GH4�R-�`�La˛r�(i��r,9�f5m:��гV�(MR��,N�N�A�X5���5OA�N��؏e$��"cF7�dt	������	P[�>�-�Z�����@s=%KɶF;|�V���ƣ�+J�u�_��ra�3�ʼ���4��$#��6�##S�l7=�j;'nxZ���8d/dй�V˰Q�+�V�t_�����}�̈6����`��e+��;�� �N$3�@d8G���[=�QmP-A����$�?���A����֟�3|o�঵�9�Q[��-���X��"��*�S�n�y�HkݑVZ��Z�暋��=hbǏ�$<�`��p��ߢ�<�Kˠ��9��U�D�#AW��T�{J� �TÖN���u�V
z��R�c��&Y�.!h\�n>1�
C�9j4�1�FWT��6<y)�u�P�+��:��+�Z�l DG��j��W��[��1ˬ�kM�]�T���\�/嶅`���bJ�>��t�j�v���6�?��e��3U�ǀ[������L�����}љx�67��nZ����2����2ߡ��*�2�bo���������{�F�ț�E�����A�\��k�H�}AZ�"l�=Dt~�����E��42�2��f����_+�8ˠr��OG����~@e@71�5��s�T��l������&�Őn���n�^����s��wLq�$?0~Y�)	��N7��GP6��� ����FPw���f:������L���{d���n,�q?Xڋ�iH���x�oA���HC�����k!G,������E����ǥ9�����ڔ���r��|<5*����l�A�#/�ʍ��c1�����Ѫ���c��|�gH.e�h ߦ�4ff/��˃�枂���{�\�K��<6����j�E A��b�C㰱�髺#V�F�w�.�ЊD<����5�#�d8~ќg�N�P�GpBd����|���&�<��
�^�O��d���{�l�iL�K}"?��n���X�� ������M42D ӈ��5$�R���n4� ��q��<o�AsC��GP��a@mX�},Ç����!����h�n��N-����5/v9Z��U~k�c�d0���d6x^��A�=���+��6�O[<!�G�J�&���2k��QJǔ�_՟o�Y��A���S��;�Q��r	  ?���jI���[�0ZĈ���'ks`�q�䣧MC���;"�Ў���,�1��;v��d�lUJe	3��+�Fj��oD�H|ӕ��7@�_J@��A�&U N]-ݩ/DJRjZq˵G�8Na�sjR�ry-�h�	����jƨ)�b��/�S!�Q�,���w%��/�U���F��v��h�Y�c&o�����%�y|�r0-L��}p/ڵ�%���$����^�Q�O(1/� ����h/z��b3�pT�1 G���EmW�ꒂ�X��Y ��5�}�Mǁ��4���{u�c�
bE㴞�ڶ�
zF���8��;�t�@��A�/;�nz#+^��_q�m?%۴�s�=��K++*-�S�g������+	�J �$IB�o��h�=o�p4���g6�'@BlM��L�� 9g��ܿ�AP}�=M%�Q8�K|Y0��O����4��߆���A�XoU�w÷@T��ޫ�,���j��@��0��搜�<�$���G1�	6Kn�V���WK7zt�zB=ۮ)o�b�- �V��L8Y�'�ӊJ>�ޘ���A�����0/-(�U��"�FvMO������8EM���c���'�kr�B�q̛�1CB�m��nd�h��C������0���I�?�`�`�2Xs#�Y�vȹ��?q�R����z�v��T)v�kI<����3�9��(���M�4�������S�X�����C�m#T�yU:F��S�x/=Q��ktm�ٙ�mM<� �	��J�ؙ�(m�S����*Y+I�����;vD�#U0�53������Ut6��������3}jN�ʢ}����G�'�ʃ�!�o_j�Yf��J���̈�|!>%@�L�⃜ކ���E� �P�m��e%g�i���$��K[�`�4��q�Bo���7I�5�b��1���Y�K���9c�#��o�|���M�<q�5��UU�����-�A��`��HqY��ܴ���V��6礳���:�Y�<[����o��C����> �H=7�Y��Q�?6u'��Aح����?�.�7���gx9�BFڍ	酊��3�J��+ �S%�+��b�4g1��,��$�՞A���P�ؗ�������6����8~:�}y"z�Ӏ����݅�L	�)(��������i଑�Z�b���ʹ��G���y�W�4zp>���57�6�Ls�ȴW�����kB]�0�4jgH\/U�a�#��q�J1_|�G�u�&V���b�V���y;��JD�S+��.��`H����*%Z(�z΃z�
�ˣl#����~<�|�չ�L�t�Ps#�g��1�O�ӓ�XQ@�N��4�gmc8���(���/�S�=���b�EC@��8M�K)0�O탨kAVϛ�T|.��������zO2/p�e1�}�6H�̱�����Y��P�qu"���I^6g���t�j��RثYvs��^Ix��t�A5,\b1���񑫰��6�!=�{#����,o0��-q���h�+!D2>l�Q"���B�ˢ�l*��nݪΘC�t?u�(��~s��@�������,�>."x�ʤkDi�P:ȁ�m��e���Q��!_`�N�k7�t�ީ{���RR���ؼN��Ƃui��Y�%�ڀ�t�`�\}j�.Ϩ���X�cG�c@���Rk�f�=����Qãc��[T0�8{O��c=���[����x�p���g�������h6�d�Ʈ$;���v"�G�[_ll��+�~VΊ��S8�_�>�OJ�l�+|{Bh�O��o�ޢ�A]^eҗ��5T��\��t����pDm��@tf\ t��u_L�ۗ��Ź�|�е\�^ߑ�[P���A��C�p���p����t��� K�5�k����"=�c?�y��W9�IQg��.#]!��l>]+ާ
�\>ЬE�J�� ?H��ܺ`�t�<(I�X�&p�FA��f���~�!�<���FG��~�K��eݽ���WZ|I��Y]Ӌ�z�3;Kzɬ\ZRŦ�m���2 ��s[u�t3.�L��L�������ŗ�8�߮�隵���EQ���q��5)�JzԺL����`���9��[�s����6�;4B6�3��)|����S��l�t�NX�Ha���[@��6%���J��J$��,�ғX�}�6��0xi��WO&�!?�}�L��L��H�D��U��ń�0c�9ߓ��3ҙl�[���K>)⚡ɦvSAN�������jy�E���*��ez���!���������ʥs�T�­�X$*�1WpWc��w�,h�A8�H B� ��P6��p�I[:��9y��"�(|~(̅�)n�Q�׊ܸm��p*�3!7a���N@>	��]? j�s7�F���O��-U;�\`-��V�*a{�n��I�d��]`'�:;��fd�?H��b�R`%}Y��^�6���!J�9,�*_ukӥ�8-����mf�[W1���}����%���8t��Z�f��(U�I5��['�_����חr����(�"������T�N��k�d�g	��w�`�a����~q�}�d�HR�4B)ը�h�K��c��]���PT��|AV���W��V��G�S�R{�k�8iM�&�S�YGA�䙵�j�W�Vh��n<�:�)�h�L5 �"�?xg��.F�O���P��}֚� �c,�&�+�G~ɢe3�-�edZg/��`~�N��X�ki���M�uC��]�/d�k 2iǑ��T`��Iƚ�1��l����ca��V�ߴ^�a{EN�H:����#�!;ʏ���ixl>g�y�+�Ewz�,2"��#Y�E�fUw����Q�h��+�<�^��ۜ�&�7�#d�c����
:,�X�n!��4����pG��=a��K�#�;B���F���c7��	�^��6�]?��Y#3N�쬬jy4��]L�nv�����g~D�a�jC�^��W7@Ii���I����}�q|r*��
P��Suy�.�Vhb�SE���_��a�Gδ�o��Xr��<�[i�v�0A�qu|~�z�X�A�I���ϝp߈�����YJ)�)����"@������Px �{2A^�,�D��,�
�q�&z򰗞3@�A+�&{jB�&bm�[����޸$�u��4k��.�^,�������a�n�$�p�ϯ���"r�/`��X�y2錵�g�?��w��|��/��ȳk�V�Z��H`���Ȭ��[%9f;r��T��r7fZl.���H�}�Ah
!-��/X�Jg.��i���'�ڽF�s�p_�Ím�6+�!.���������s)�t���@јE�M���+�hQ%�=�}�62AD����� �`px樒.��E/�LE`u���8ӳr�oY����m˒YM�o#mj����VYk�;�@	���xR�֟�J�__l3*b/>�����-��zO��>RF8�� AgE�J%~���Uh�g��u�A��`5�ag�w��L���v?-ާ����q��� ��)����-�����.�ܿ����=P��I�O�
�����j�����w�{6�U��Ƨ.0�t�_D�h(?�oB���%>	�a��f� *��t��b��1�Gt�Lٝ��N �I����j���H�51��Ml��Wf)�c��rL��Qj�Γ����'�w�lf73K�k���I֭�7N�7��iF��4���Xn.�~�VxEJ�Ԫw��_��U��ʀͥ\I'٠gCw��d�2�7f��ƌ��F��V��{Y������^����Tg��p�߅� -��d�7x�������lI2�1��S�y����U��ꆎ�K�2@�����Y�(`�$9^1!e	��`hssN=�{S�5���j	����G�M��)޶e�J�F��I���O�R��(��YKg�JEb�GH���9�k������� �-��%�e���ӳ��
Wu{*��-ŰO�z��� ��X��mrU�����+�����oNL�fa��P�i��$6Bs4�r�̓)�m1�'7VO�PL/P������/
�̍N���Su7iܟ��x�7�?:4Oߨ2�\aq��-���Y9�<�Y"��`S���F�Y���))j�z��sZ+�`BUKDF9P8����
b)����n_�nT�0>ڌ����x�6�bH�Y�A���Č˷����!�Z����m���0�����K�:V &
)Vh#�9ӹ��1p��i��NF����J"�BY��Is�{ن�1'{K���c�"�N����%�<�"�]ǰ���P彑]��y�	�eF�Xm�M����k��a���J(�_G.�l݀�e)=�J�C��A�J��lA�}&��l)�&"���{�DEq��x�t��Sk%�l7������Ԟ�F6�_��!�B�gh̍��A����Z$q��@���g���S���MG���n���mE^9������)�S���ضr�`#-��uc��3/�"�urv�4�5Oզ�n���/:
�O1 I��
�T�"ѩ*Yp��O?ߵ��wy��ʟ���ɺ`FXR��z�J.2"�%��ɍ8ؽ�z�{@h@]ǸH�$��u�ʧ�|����ր�Y�T^��CK��al}a����@Y4}�_w�l)�s��M�RC�헜%J�����QUZ��98�U��e�Z�Xe�8��?����-�&�5�ĩ�/Uذ��Iteh}����h8�&�sE��� 	�Z�z��ʐ�U��	!{�4�ZC�.�K���QaA�|+�p���~��k��A�S�ุr���F*��vS�|��(c�^@ys��[��O�U^�3C��)R���a>����"�G�Xo;�'��gs�~p@:wy���ܼ[�m��?�{�������,e�����q�j��:�Q@�S/}Y���RG�������R�Ǝ3r��W�|r� �D�z=�GW��Nq�@YZ���fwd�Q�?HH-
�����`��ݕ7:��T����df��g�V��DA�O NA�՞����(��5r1��~��\%^}۹���m�~��8���zÂyK�I]��в����M���*~m4n�K(�c��T����Ý�O�c��KE�(j��Ktg��w��J�|%W.)f���566X
����2<#�$=T p􈝳Q���/� ����2�����Z���<n�*�X�5����ƛK4�g����ˋ]�����1�q�(��[�����Z>�A�8Ѝ0�S�t�/bH���9����=m7U�y��!����g"��ju��H;�;%���H�b�&���~`��}i#v�D���	�c2$�ψ�l�E_�`�	�`��1�np� 2rOP	����5�s��������V�i��W74�6�Ƥ���-�'4x�����"V*�̞�������*,�)�ڝ�e��j\�Qy���?�+�?(�1�]ݧ�5����/8��G�����y�����=ت�mm�M�B
��/I�Z�@&�G��f�V5���.+Bl$��6�&%�+� �H��G:���?k�I+M�*�=ynq�L�a�����tw>�j�B�Y�Y�O��*�}�������4[E�u��.F����ï���A=���[�W\��������`�Ǿp�ا�3z��-K>Ml0��̂jQU���䯛��DȢQ����.��w� ;J��5��_�Vx��ik��U�A6��j=+6����d����/v���zTZR��t� i�]���{~Q���`�ϋ�:{�v�i�)�^c���w.��'���Ŷ��/�o�F�.iN8��*z�<c+�]�rէ؊��$N7T�8�D����@|�!o���ݖ����A���z*h^i�����>.�v�.��e��=cvՇAY�.K�Η�Q�6�	�w��ɰ�y�ub��8�0��x>�[6�e�������9��h{d�N%����@��Ų����j�T�j,V>?�ϯ_v&�؁��m!�cW�{��ہEc������.�Nr['���-m���Hi�&9?����FiwK��2��\cj�O��k��X��h�|o9y�8C�i^���,q_���r��w�ə%�=�S&����H��ߍ��A?p�����N��e`TM����ɥ�}T[Nv��cR�K���@Q����q㢝[�H?e�^��j�!����/��M�2&$�G���n��]ݕ;�bP��9��X�KG���}�]�&\��ְpm����E���|����#�W��@��Q}�;��&�A�8���Q�1п�v����Pw�A�s�Lj�ɾ(�IP5?�[|Н�9������l��o/!:�#��95���p����N�)�,�\������kk�C��}��G�֞h	q��a�
sȁ"��
yn��I�,e��2��C��_~�����^�	}���Q��gH|����T7��K�J	FO%���%u�t�#��C���-�\?c���Z-�I��6�ؒ]�b@�O���a!Q������������҄�ʫ��a�O
5�rB��Q;�d���J��=����{gw��b���P�,&z�6�SÑ�����g�<<^���ZB�M`l�e�1h![!���Ň��ՠ	�3�*	��C7�%��'R��L�/Z�W��~~u�K9�yU��5�v��ț��M����\����Ƈ���	q]p�x��|T�:1@;lN��5!C(ES�+u��"� ��s�,��	1����%�^ts�p ~��~!����~(,l��wa�NM�dQ�z}@��yvk�nl~`�ڮ�6sj�)a��M	ݿ�{&�Ι�^A�O��;��o ��6����lc_�}���M�k������V�B�w�Y�4�$m�` ʨkg�� ~��<t�l�k��o�v�܃����R�ܸ�y�d��A�U(n�!� [��d[ ���fI����ō��E �Zd�LM�/�h���G#�˥���/���w�{(p8_@��E��',6J���A{v�r����.B;F�ymOAq�d�x�j��}��ךM�B%�PG�4g>j!�=��hw�u�i�AG�+����ߪm߶��	�����⩆ӆ;�d(z�3%���
Zu�1�B�5��������]�]��t��#�2f�Ak��^e���t�K��E{����&L\�Ev�~�V�1��GEC�x���q�r�Zڤ�W����C������K�565D!O���M��E�m�,Rh�3�(�E=>�������b�ڌ�?�$y��g�R{�|�}9�ʃ`|�iK�w���H�hF�5Tz���&�j�fa�u�Fṁ�I{:���^Բ���L�\����g,ɣ���v��ài�ln^E����=�XZ$3�k����U����e�@;��P`!���	�����y-�+a�)�,�ȏ�'W{��>͑���C7�H�<;1�o�v���S�.�l��'�+D�����Sv3`�&������i�q��&7�M���%2��&�\�����'4s�{��x���"8�9��Ϳ�$�<�Y�A�~&�dU��?u>���ce��ؔR�����,�y�m�C�,�9�x����I|�kK��.�n���yW��'�NLeEV�q�l/���|�#�IQ<S����V 1/)�>!,	�Q��x��Y6����afR_��FN(��^ht�x�H��?�ȱ2e�f���&��x�s�CR��˸�Z6E'�=c^���W\�þ]q`z��]佛���7�s4@�ү������б��+Y�t%>E����@�v�Zp�z8	��t��K{�sw�{���q�5(�n닼�iuS�M���l �k����U��H��:_��{�/��ߦ��\�U�}L�hO����� -����{Ź��x)S4�(X�eZT�!2�� �_3��CZp����ظ!�ܸ�+f�zdJ���b˞|ow"�u�*ót2/t��i)5�߿�x�u��x�����~Q��p�`Ҿ4n�E�7B_]��db���h�1Ů�捾��] I�ɿ�T���*�fCQ��nR-,"\�%�C������c3O�}��jG�� �MD�o����6��<����D��**��Sf��îccp\c�f�d��+y���� /��9lz��@
��'$q�8�'��f�NN(�r��#��`��9+��v�������ۭ*�9c܈�콭3� �|�n�b�](v���8�Sv��6���C�o�� L���[7oE@GRK����"B��T{P��qi����S�&~b�}bǏ���}´����� ��d�A8���<�������'e�Zow\�,�<^�B�)���T��ƀ�p'����Xob�r����O{yC	ID��M(���3w��H�*�����ĝ�'����y#!�/����n	���`���e8:;�w^���SVh��aoL�U��vP���b�pd&�BD;���U�gQsJ۴S��t�x�2�yF�9-��� -bz���DM�s]?�- U��(���� AN�o�3� �ɕ ���H���q�.�e!��)��& �G��
��癷O*;��ېdp��ٹ��X�֋}�0���|84�v�F'
��$ZtYA��?�W�v�`�?�o��Z�k�u���U�Ŷ�:���6Bm[w���՝��۔��D��:���� �/n�*� �:�$[eF��~Hb"�+ ���{%+�A<!�tF~�5�NȃP��y�8Tt/�&Am�����k|uC�� ul���2���ٞ���*���?D��r�	Nd�x16�n�i��Q�c�{��C����%�F��aֶy-i��ܼ��ޜ�`��}���y�p=}4$덩R*(È��`+p6{j����	��p�A�d���� �)c�Or�73�Жm+�'��#� ��>'������K6�9A#�栏'�Z�s&�Vv��Kɲ��Ζw1�Hw��P�F^Jѱ9�����r����V[���m���a3AV�����2d��"���q�#���|,��^$�s�Ϛ��܈gI�KyC锻mҼh���
"�%ฉn�Z�҄8�j� �ꮊDd&��iL����[
�;��%��'�U�S.$�uG�m�����{QءX��|%9wU��}Pcԃ�@WF09f��<�� �K���~ҿ�"뛼d�4���[�I&q�J,�-��ϳ����_� M�L�q���	-֍L���/�$��	]��EvÀZ���]N�Ȗ��# ��|����)H����������&�*\<���E���[������/��2+��r���2���i���/yl��5|�W+�BH+�P�e�9�#��c~*ސ��:n�,6����Ɉ�Q#���]QJ�~W�xs�5ݨ�V�J�o/:���OlLq5�*��7m?�Q�N�9B�,K";|H����$x�8" �͌�/!�=^eL��<���i���$8 U*����1����Ƕ��kߚh٣��s�2�zo�V����tU���	X�Jn��M-��  �J�p��J�E�\+�Q٦���c^&��\3���b�~g�����a�?{T����G�ܹ�CsT[�f8�+N Ҍ���2���_ڳ�G�b�k8�N������G��V�}�o�Bͣ���F��Ҿ��ϛ�X�K�b��	�0��
d���E�*�0`?���wk�F~��I�;��W)A%�ar3����6��7���>�X��g'�K?��w�b�]���zQDM[]RHm
r���7hs�-�j��X�e�xЅO�U���X�.��ý��׾EHM�R��8�{'<�k+i%�d�rr�d�Ex9�E�֛���S66��)�K�ݜ_�x
��e�CK���V�u��zR�9U+�H�!�ќ��h�{��݄��FKS+�du�Q;WF	��H
�F}���5�q�!ӄnz4��@�\��a�Iܪ���$��慎��κ�_s�V^��fǑ���:�֬S��h�#a!����6��R�x_����Λ�2{epB���]�7�X#ö��HJ��Ҿ���c,���2K�����w�(c�!@s!�4�&H�^�"Q(���������z��Y�`z�D_���^9���?��K�w	Z;y�Pr�D���8�3��f�P��׹��pݏ��ǌߗ�c�c����z�PS�l��6��f����G����z6�l��Hl�Sɴ}�؞!�ilO �/!�(Q���iߟ����ƕ���1�g3C��1$fH�uأ/m&4�Ic�G�0�Q!�"ǸM��F�P"���Т^�+a�1}��H���(���D�y���	Jyv��!��î���@f4*|�I<�`՟�MYO������6U��Ɖ��
 �f�1���ʔ�"��Y�.6)=��[��\��kk4Q��lp)�)���LHk)�X���$��Ќ���^҉��sU~�J�����k��y�x������\� 7j~۫IUuI�~Ԃ.�x�Ԏ}Έ�'O�������*`�l}{Ѹ/� )�_D����6����6��� ���J��֮�ui�oZ����e�8�؊�d����uL���4��<�'��<j+��]�����3�-;Y{��wC%D9�:˒�t���?ϵk L��إ�R(f�Ly�%����Ӡ���2�Ye�f��I+S
ӷ�v���Y%n�j�۞��۳���D�Ή�ݔ�KM��p ����2������1Cy���"���W`^#^��P&���ƫ�Rӓ�������
��9���9����C�[����M��r{
�X��W�@^.-�_��ֺ|�lle�+�<	%���S/�w9w�E�f]%�.̠� .�p�iߚ��*}�r�V�����=$۾�k������_t�v�H�3����q����a�Xg��V0j�[1�ϓV�j��	0KAYt�D<k�ֽ�2vf�3&��;�rq��웪I �@WY}�ۙ��#}��x��W�Q����7᜝Վ�M��/)q�2��B?�Kz/`!���С���/��I��V@-�� ّ���F�)���ޥ�\#5������ #'����&�?���4_3��~I��)[�q�*{�RD�S+[�Iu���Q1���C����w���^��Uj���6*�X,f1�rGc"�eCC��� ��r���J�;���dȘ#W�6���yh�@�?�_v��?~�Ш�S�K��l[
��&[>�:��s�
��N����9~�3�g�N%�=l��'%--��H�n�E)v��u�:��uW~r�ʒ҈��0���`�!;�y)�L�S��L�T�h�����(�ˎ��2?�D��RP��v����$���_����7p渠�`��� �2�s���H�S��H#o2�n` 3(��N �Ӥ�R�-��f�2 5Ş4�ze���q���Z�0��Gupd_(�=)؃��a�R��WBM=[�?y�oj��sZ�ᓚ)*1W@K02>
ķ%Ӌp�Iv�(A& y{��}LFVDeI[TgMS����h���=���ml�:����f��ͯXkb��-�R�{�%<��{h��������eww�+`� �1�����Ge(�<�cy]�3����^��f%�K�^��b��8���-� ᕃ��J�>x}��aC`]�B�v�JI�)N�A�E4������;�Zoh�;Eջ�K��,��|+<S��r�~�}ԍ�����_������\�_9}��L������Ur����C�sF7$��Å瓍���s�.�:n'��"m�TF��of}���V$a�]�騋?u����V#b�#�>���Z x:��c�'pޤ��cK9�O��愨#��`�����egcl� �^8B��@���ࡗY�n�Y��I�TW����Сi©=������<�J���W�U�&j|�Q\�R�,x���.Í�9�����?�U�ښW!�$B^7��o���v����Z���Iz�r�d�!��E+E1�\N^��N��)3�O���|^mP�a�[�ݍ������vX
p��O>�  �s9����"
<'5׶Ru��t�(j%�/v����FnA{;۠&�'c�8�A?��*5��M&�z���Q�e�<q`��K(r[���=]��kk�x�A3�P�
�]��ҕ�fƥ/9�����厳1]�> ]���o?K�-�/�nI|�횊&f�3�N�x��z$o5�)�gj[#��mB^�B@��$�O'Qwk���ҒqT�[�y|��WpdA� l�S�� �✚��k]�>����'�L�qˡ�^*(��K1��n�W_7��E����S-L���+�u�'v���~�w��_�՜;��߉ܨ�F��yC�9��Y�a`����i�9�q��&Ǡz�U�� ��p�-XG��q��iJ�娪�B/�P:�&>8P/�M��~��P�S��7�Q��\ح�4��k�7v^�Í��5�}�f�t~	�T��b]rjC�53i�`�ϝ����'�ێ��E�8L�լDM�
�Q$x�4���j7O��	�z�]��;�lIG)��,�V,����E߅k���D^(,8S+�KI�CCTWE"30�E�*�P�V�g���\#�5z���_��H�@N��g�J�7�0Gߴ笧����b��ޤ����޵A�<9}�RZ��R����]G>��sW�e�%�5��?��@�rO�vp�<@�
��w;�P%@
h϶��'n�0�/�[|'��h��ԑ��e�T:�w� �<�� ҩ#��qQ؈�ѕw�
w	���IAl--:A,���65��ғ��S�ܓ�1MWFqA���``>�ُEO_�C�n!�'�0g�k�o�� K�~Q>C7�x�K�sֈ�V?�|���;�w\#�P`ɲ��Svb���T�+N����C�_#Q*]*���Q~��X������)>-\]E�{�)&}W���S�Z��Kᴙ[f���d:�����W�%?;�⧙ѐ�P����c��ik�v��Ytu�vB$G�<>��iZ���M�҆��H1��)��ĸQ���Q9�� @�Z���r��P\�����[�V��6ZX��	u�)[E_�Y{�}�䴮�}_�$�̼ �k����6t�6�(���\�
�	�,D�;1�&�V]AMSc�b�����[�c1[��ʳ���b�}��)����f�9q�~O��,I�e��;*DI��^� ��/���x���x��+ڏ!��/qUc��f�����#��!���/�����`(Ip����I%F�v�{�w-���:T���0�p}Ju��.l43��,^L�eYr������/x��W����=��>^9m���z�|�ފP�&~V�.�Ab3�X��a���Ǩ�VO_�Q�j��R0C$z�s��X��nOM�A��,�����s�p�1����?ݟ%y���5��A�
A �r�4��h{��m�T�T�?�Ίߘ��q�J�X��~�ԓa[#�o�[$F�����c�}%��+�� �	XIX��lH�'0��@�a��8:�5�����$}���,Huc����j�3%
�@��Y�Q��f����3GGu�B��Hx\����iOud��ac�H�H�f�(>C�U�?_�����:%��o���It;~馲:G��:����HK-�%+��pkj�B�7��g%�\v|�.b�t����o⟖�'���	��q���ȡ�OS�X���x�[Ԁ4�YLa�"BC)i�gԚ���̻Rc��U(��V�z�9s ���[�U���$;�.�Ua�K�w:��9t0�TPQAzx&!+z6��vh�:T��(� ���T��O��N�7hP<>�������CS�P��y�p??%8Fl!4.��.�F�$ͩ�)6�2)<��a����T�{�ѣ�1GD8ɩ�lF+bgS)6�0�;0���-����r;�Bc_v����$���"U��y�q=LK��,L�Z`�H��Y�Y4K��lNF	�y�Fe�� q��4�^Y���:(�T���K}ǋ�
����W�h#"���Bm@�E��6wA���ӓ���(?�o؊��,̩c����;����/�<��ɑl�D�9l����k�%�|�Im�������-T�����J�����L]����K��Bѧ���.Cy����`��SU�@_C5�L�cO^����Մ�����#dݺY0P�X|�?�ܻa��7!���wSaɌW󘫢�*�	"�ڏ�t���VEf�M4B��
wsz6߅N"�J�5��=c꺒����&N���(r�9�$�-��
 �5"��Hx�2��FtW�����	�|:�F�'J[-As�z�����9Eݓ��UT�C����Ix�;����Z��0\ 1L/g���R��p k�������2P�dK&�8��I����*A����K]�a�������M�M�g��[��<��%�G�6�ʖ|WFР���dɐ��7*�Q�騝)q�H�TE�d���:5�h0��_�y��JQ�M�{b��Uں�ˁ��p��&��(����ë�����*p��<�
� Ur�5��*L�-o�T�� `[B#e���f����.D�.��z����;��7���_�O�H�o8$�v탨�]�Mwdj�։i�|���`����y*�?L���i��V`}E��}5���O>x�t�޻Ť��W�ﳵf�0�'�ҫP�A�l��.�~U����@�w*غ��!��7��f��cI���<�ʐ���ء�[ ��Ksݙ��ܸ�]�fe��ߓsU�'��>�/�:zG��w�u	ns��Lf���{�v�x]�?q�#�6�p*�Sm2x�p�>�MEj���t�#V��f*4A�6xW�3gX���L�N0OEˊ��l�@�K�܏��	�n�����+�R�py�*�r�>ώ:�GeC2Ê�=�w���u�^
NE�th�(%w�J<���ŧ�qگ�p/�EB���Y�$=��m���>�W�\�I�����6���,�����7��G�Z,��3��S��.�g*�ch��d&�O9�9 "��r'R^x���Q���
Y��	PC�Is��L��U�]��s��"Y!U(d��-L��n�O&t����/�q�t�B�����Z��݂\��aG"���J�&�RA�,G������1N��Q�d��d�.�ҧ�ı���#:��i�rx��e}�!���0�|\B�N���-���y͒��ۙ}�`�	��H0$�<0�d:�0@��Ȥ�nō9"�u��28!|��a����P���2VA�f<�GE�þ�U��P�s��_�&)0C���4푬�'�L���
��#śR�R�I[(���tu��#)`�~Z�I1��=�}�a*�ƞ���|�OS�,�V�m؋񞂹�֯�������[�	���� ��'�L,���8��p4�p5qm-�,9�3�_}�H�!��9����|�O60�^������-A$�wGR�j~�ɺM=�p�N���h�󾹨���r�'�1B�1�,��4b3��8Zl�� @&iN�
e���7���h��#*U�4<�?�3�0B��M���^i(�rsR!�0�&���S�?H���|�h�ߔ<y�w�Ι[�}����O<kj��FG&a5����K��G�<q���گ���ߋL��gCD�f��
-$P��?�fqcF'��v�O-��u�z�+�&��Q7�,#��Y��\��Y$��>ږП�ӝ�s���g�,�:�O#h-�^Ǵ�D�9 ;~Q�}���6����P�p7�P`��?�ǫ�m��M"n��cFO��aʹw%vD��Ҫī��1.��^�b�O^@+<������L�<���dF�"�/���%d��o0�.e���C:�M��*�8�c.�̟��ΐ�Oі���1��[dJ��JVwms�9axp��4νH �IZ�a>���0&���8p-[JV!7K�r]r�%,�Yv#e�bF![�
i+辢@Q�()orgN�N�ڏ�����g��+}��|�$�U�"֧�FIBQ��7�l\5gd�[zF�3F���g�,ڷ�o��X7�{$�u���]qY�O<�&M�D��g���g��2����������^���3�Q�$��9�Z���ר��6�vJ��,���:�K 8�a@&�[T���ߐ��U)G��T��7{ d2U�Y�"�t�f�c���@���[=�W�X1��$�*����mJ�a��)g�����Vֶ���gB���QX�,[a��K_:蟳>�SjG�D����kIq��)e���������Zg�(ؘ�x~E�z�����ߑ��q�D���h����W���fjs��j�3�d�����g?��(���h�HuA�\s��o�ٱ�?ͫ��W2����������+)���2���D�EF[�vU���d���;��,T�Շ	å�)�d/s�eۗ?V/�>���W��*�eqö
���+�A�u�%o�VN;wb���˒�����'�?K.�|?s"������k��s��.��y��?�~������.b31�4�tl��_ɉW�`�����;-���t���y=U��ޝ-(��DszU��׸���-�5�t��h�2n7�a�$�:H��:p���2*�ǭ��fwnۋ:G9ju�s[B+٤��#mt�R�jY�GwDh�@�*k�N���󆺑�Τyq&8��Vj�l��ҏ%Gw��x�BX
D¦��@-�"��$���<����j#�G���;RYH��%�u��U' 6�)��%��{�\�����0��r�	ny5�w��m�J��K13�<��=�.$�h�H4��"ˆ�k�bf��gh��z��0� �>�y��&z����?.�-棆�D�~�V��dHZY��e��(��~���7�bԪ��Z�ڱ~�'��4:h?����Gn�ʔd�I�<���;���������,�.F_Y:��a*���(b!������;�a��4����ؒ�(��?f��(C4�Mphș�����ZP'NE���
��
TgN�[Y=�j�s~���h!V��H���"�id�3&��Z��v]��tn��6�6k����ɝ L��%g l��[>��S$�rP7���ߚ+�������k���ʻ�$�
��y�7���6QgP5���"��rq~�D��RՠM�j����y���a^񹐧8����SZ��[�ll���af�n̝K0�_�ԗU��;��3���|+	�Ⱥ|�"5��\�����Z�J�d�#�}����I��=��f]�#�=8C�b5\�Z�M��|����
OT�H�[.����b��i;�]Mf�1���L���Fl@��kԂts!�G��حG�17��i	�=F=�'o�9�	f����+��F�A��(�� 1Z>@���˯^db#���d��܏ሑ�o��.��9)綣���(��5Н� ƛb�d����<=�	�9�n�yQ����.��ч�F�Q1&�T��i-"�����ˑ��p ����Qx��v�]Dr���|�n�F�D��(�O���5b��\���W��r�`S�6���t M��K�>/]��q�m~x�+�Z C��rX[bn�4���t�U��T<g^�j��xx�FȡO���u�a�M�_쾘���/�[C����Wf�?���%F�q�FS��]]C����g���FsyV�/���/�YYC1`f�_D�{3�J�\u[}�'^�rut��!��r����o�r��U���7��kZ��u�I���.��\d�E��֖�X�w�%z��!�l~�=0�
�\fp�Ht�����X[5H���Y�Ju��01{叩E?��á�>�����s:(-�����y�pƹ�W����8/���Ц�$ت(+<�����?�k���� J�����@�8�5����2��)��ZFUEר6���jj����h6ܱz+���"��2u)��<���pRſ�U
;a���ݑ��\Y��`E���r�>s��{���e�-��U�|�{��+��kޜڗ� ʫ�:���k�4���ŀ*تw�'61�p3�ZQ)�Sx��?�����$���%�n�X�ȗ[u��l�AB4�t� �-�Ӎ�L��w0_u�>L���g���}��n�hڻL7I�N��Q~y�����e�ڠHTih�Ӎ�H9������z���u�{{U�n�>h�f+P�0=��>d��r��oUl�$i���fh>�i�¡���f��,�eQӔ�68��D�^��mR�t��).���v��Q�x��u�}�+\�{CtZ���VD�7љx����&A�^k �Z� 9RW��Qڠ���Th�< ��RL�O��y�;�כڝD��V�xʛ_w�d�]Z9ZY�+�rU�#�vm�E&	\ϡB��Hri�9&~��+���ҩ	S{ݷ5�rݮ�8�jm]��b��~��$T?Of�)������߹�Q��N�9a)�b��}��~���A���	u4Y1}�1��)K��EBjk&k+W.~��H߆z�MN�D~j�ȡ	��O>E�@�_rFY+fH�����m'�o�gi�E�q^�#���@�]~8�:�/��������ֹo�=���q1�vM�w�@P��$0<��p�PK��v��#`.է���
�,�_�'�w��������Ѿ[R?\n��]���͢K���H����2�#)�c��8�m�ۺ~�[(?u��U��H�Y]�V5�\?>[��A�iW'�*��5���5���N�O�@��,�YY2�Lm0�+#oØ��"AT�m[�[�"�ZܓS���ġ�����|��N:�v�U����'}��Gu^B(�a@�;�-7_9!�f�U�]��c� �D�I4�� �^.��6��\'|{�����N�ibEߛe�ɩ:�5��t�@���w'6�+�V��'��"H9ݲ��^£�ܳO��_~E��S�����������^<��#��B`��S�6�ކV9�8Ԡ�_�(���$��I?�~���f�ܨ�0������:�Vc�~89��N�4Z�\|%�a�G�wD�6npgŽ���L$�;�)S��.����[3�x���m�#?-���{��W�+PwZ�WiF17W8�(z%���� �6��]t43�W��$kX:���^�ݩ�����.#���h��Si/����k���AX��8@'�Y0k*��^�[*z���ݾ�����ֻ��,NDH��RH�����ܤ�Fc&l��Ŋ;mFB��J ��&�5���͝�N����bF�0��^n�M�) ��6��⥱�O�v<��B�Tf
��CZ���
�S���e�z5��8]\Pl_�v}!���j��# ���$�2fK�y/�;/��z�V�K�Ka�[d[CӋ���6�j�����h\#���1)�?g��W��X��`�)�����^��S�B,]>AZ�t�4�+S��+Ꮔ
H���aD��T K���AKR��5�@xD*�I\�[�G�4��~�3����;�!���AR[0�p�ƶ`�MFZ�fe�� �����>J_�"f�G[ ��/09�R��z��GX{�~��_����a��vl�h��5�Y*�X&�~�`hp^k�6Ə�v����ӭ�/5av �]ä�?�_�0p��y����wȎ^4g;"3B���Jaf��AFW6�_�	����5�v�5EW�gK�p�w(��Q� :��cN�	��jEQ��l9�D?�{��$�C�l��YN��j������#���֍�kY\Na���N�O�JNW<�9��rw�_����V�O�
����=���Y;��:$"c�0��>X%��j}͹�Y�Ev��ya/���3��!�l��$Oq�,E$h���A���5D}�U,�F��;��(%|�ɮ�o]��W&��J�C��dY�m��Wj)�q�. %�C�i_|^��-�Oꮜ4��x0Q��kfy���rN�}Y4ߍRO����!C��K���$YQ�����3�0�
 �>��+x��
�_uЕ���y�vK��⽿^��͛�OV��w��˝6͟�ޝ�m��f�zXu��L=Ao|�1�8CIT���=y��x����!��名�c�y��b��0��=N�s�i������S��� ��F���Ԯ;e�Z8��8��'���[.	��5=��O(�k����ZR������e Zp�p��!I%G�[��?�����6�xm^����!�bB�5ݎ។����m�]�9-���x��"�0"��ֶ
�~��ސZP�ؖ�d�E���.�i��!�S�9w�dHE�\�d���Y
�l�5Ǽ��t���2��v�#E$z)��
�ǰ�Qk3�a��7��A�f���rS50�=z��)%)����i+�l`>�  Y�Ï����R�ԃ�{��r-�ΟA<�N�		Re����Q�$͆��Qɉ�>+'ć$�B:��D����A�yt��
5��|e#_g1P�pE�~�ߦ9�@-�.l�V&#�rQx��iRA�qfF>1<��ykR;�S	������g?�R2y��In-vI)���u�����%� a=��,7�%�L�Z\�Ɂ$���9ʌ�:"���Se?4���0P�x��#0���0���v��x�G�5BC�U
�Og�_��fԉ�E��HVw�����ׯ4P�Z"_�:ꔲ8��SE���)��:���X��6��ï5ه�$|���px:$[PO����q�ȣknLI!d�����d�.Л�����1v#{�qph2g�,A��HXWʑ�SN4���$h���l�·,@#�^E�z��TT�3��3�ܕ�(���������������w5����	��� ��/1Q^R1����{�[ �zۋGZNZIK0�:��P�&_�lGg�IG�����6�3F�n��~(ky��?�����`�V���]�PNu$���j�]�]4��Kεy��,"����Gʾ�]�{��ec��v5���
��Vݾܥi�[�W��w���?�������%�99��;I�\���s�ؒ�m��� R��bS�4�{	��68�ڟ�{�:���U�Q9�������+�
�,�M����R{U8*DJS>����,�"�A�/k�uiO��0}�R�H^�K>j�gKv�� P��ߺk[}��\I�|����9��i�I�Q(�s��PA��F���͝���"6��E�������ʢ����v;"��?��,�cz��0��5'�ݓH!=���7�e����9��:�c�~�]�}쉙�B�j4�K���O���1w� ��P���?�j'�!F�_.�LjX.�����.��e<�ϵjϫU�?�A����w�pge�Jx���͗����i��S�f$�+�N���������,Hk/�Qa�o���6���
��d�]<��8�� N�t}=���~��5o���H�f�����c�K�R��o�_TC�.�%	�c(\��J2} I��H��v���7���:7WRyf�Yo�t8Y=/*y�0��H�HB?��� ��i#� !%I�K�����?`�M{Dr*�^L��k9�D��.y�	�^�<�ι�HH�k@w�&<�	��N+ty�=�{�?�0K)���D�7�b���`4��5q0U0*��J֜�ߌr1��N&;�hp;����2�2&�1��7)��W�w}� ��G���t�����[�����_���>ֈ����a����=/4![P����\�	&��"��I�F�bDVr4���	 ��"b�Tަ�D	�k|ە	�i$Q�i?��
j) ��rJ�S5 @↉)����LM%����\H�^r����{4
V�>�	'�L�˵�P)����`�棥�
p|���Ł��1�Zh�Ȧ\� t,��W0�W0�l����S���|Ҏ/) ��;���R1<t�U�?�0�A�3>���%�/C�OP8�9B;7&�B����o )r�3��60��]@����������Ÿ;�BǍlX�h��(^��O�?,�y� �Aa�p�]x^O>�!���}qig%���Z�vB���.���ࢥ�<P�a#$=j�.�b-��u#�r+��r�y��K�&1'������o���H�716W�����*VpB�TNq-i�]%�����CP�m8�T���7�;��ַ���%�!Ȋ���M����������~T@}u������F]�d�1<x����%'���O��_���<L���D��?�����k��ټ���|�N��Q>���Q<����
Ĥ� �?w�R|ʱG�zT�px��h'wx7�aܓ�sK�R�}^�˿��|�WI1�{�#]T�5����I�F�Nđ{J@`�	�uVB�X�x�h�{t�`�$GG~��*�פ<͜�����}>�?��2�9�sPUZ5&n��5�~I�"�S'��`-��5|�*D�q�]�d�s�[?�ċ�����K�B��p���0�0���A�m���ŋ���S�m���;ǁ��E@^���8l��K5�l@�P�O�m��C�GS�x�Z�r~\�#���8:�ӂ��4j֜z#�=kEۻU��vf�l-љ<?-��:�U��btՑa�1��v�_��H!�[=H,�x
�����T's�]<s�;���U���d�b�r#��8�4��*��p�F
##�Q�Z��'=�ͺ����4�a��;��TzYzǿ�zo;1��`g��������/e����/=R��M.b������CylL�HS�7�>�a�쩪Oagjz�+��0�}���$&U�ٱf���?0��0����Ѷ�74�1܊���e�-����}P��B�n�,i{��q���pcg�'I�cuJhD4ntb�1�����\�B:����A�2&�<�Z<���fP���v���O�ۛ�M#?���y�F�un���R"�b��T�Nʷd��E��Ω�|aM�?��U�-k�ضIʈ6u���^���{RD�||L�>���4�la��c�����������G6Ä��Iq�&E9���Q�r`��%�Y�L%2#_J���\������?�-՝T��PH��۰�%�_7�j`ί��~�8��3�w������?��"�9�'�	3��$_'� &���٦ć�tm��SxI�Z�)"�	(S�R���Ԏ���VO��&e��?L~�"N������tN����C#�Ӎ8m�E�u<C�-4�hlE�	΢�P�sNp�ą�Яh�~?�C���&90�N!Ԃ���ԍb����
�:x�'e�$���{��Km��,yj�l����r�I�Ud�Ft���o���n�z�$s�����2���#xjO�3��w�<Ї��Qq�#���S���jLKb�NK�B��Tn0֓U���Z)�z��4�wG�*�y�H��_�U�y��~<�d�_TI8'.a�hX���D�s|w0h`i���V����ػ�ğ��܏��s���������}��f�0J�t�4��L4��#ů� �.V\c��F�qFSr�������c.YE�St}u������Y�Z�V�q�'4���������_�Ȣ�����dx}��!$l��ry�W)�,ü���w�^�Kb�7���@�����#�WKB�^=Oia����!���g�
�f�[�� �o��e*�M��~yY�΢�9*?@�V{�/���%և��7�6���T�C��fH\��n��n�ͺ���,/�~&�i�1��[nRF���2C����W�ɫ X���)�t��<'����Pd �o� �n�ge�&
,����Eb)p�%��M��?����ز�hfbS%�J����I���G�M�����TJ�&�N�&�8l�[���, V������K2�/P٧�G8�<�HK(������$7��LF,�O#�n1dƉ��6^f�p�A#Vy�;0:">�����$��tu�^�v��*F�?4_��n����>Q���U�,�N'�ܜH���O�#��Mo1,a��4�+P��$�\�����T�.	�l-g��5@�b�I�_�W�iz�	[�ӉK�n ��r=�M��"��5��T3Z�<IF���o7ٷ�7��O�;�S(s2���f��?X�߂K��G�Mݱ%��.p�dL��%rxL�d^��8�o`�=����q�%.|  ĥNF��<e+A:���a��)�/����C	�-�3�/�x��Ë�F�������SV;��Ax�@�� ���1Ψm���+ir1��`�!���_uv��wO��[Ri��>�VD+5�Lk|[�OyTB��
��,gՎ����gbe:�}����G:�D:������P��8�t&��U���I����L�(�W7�����0S�+�}��z5|�+�L�܀���X{M^R�~�P�2o_2WLb<2*S���5&H_�`c�P�<̖w�����n~��}�|Kn}c�]H�rA5OO��W�L��D�	�w���E���<�N�m�,aS>�r�t.�~���!�=a_+�B(�zO�`�A�2i{���d��CB%'��b����5Vb���c-�D��۱6��Ar���䑔v3^ �v�\�Wt�Z���;x����NJ���O 8��+F2��7�.s����i_v"8�I��?����Ϫ��{s�@ �"=�;'��u�Y=$t��ۻ���[��l�c� �h
7B���ޭgl_��o#{�e�}9iIJD|���U�����TV�~-���hJ�'\�	s$��N�`Ƈ�����;'���&�Y@Q�R��� &?��
��}��<��S�6ѬD���LA(-��^��Y���ֆ%6��3�=N�Ā��x�jEf�#�yS��L�<1wM�a2)T�ꭏیql�H�H�dE�:�t����d��2���w�5*a;:ʞї~J��L��'��_:,J�fG��4iX@Z�G�{��\�ee%E����k!����n�
���^l����F�̔ꧏ�_��A(����U�TNk�+����y�{��&c1�;i�yЦ%H6��������"k��)� >�.:��&����������f⍊���WZ.����5>ޤ�;��+i��­��0��9��K�jE�(���[wZ�J��5�������M�veϱ���Vt�`�ep�~�ak~/�肑"�kd~� ��41�*x��ox���z;ϧ���V>��c���l|DS���XD��Y�. �6,�hvB����� 7��1�W��b�㉿O��Zh���?54f�,�hR�Ա��|t��Bچ�݊K��i*����B�#�m�k�z���m�Q�c$����3Q��1Y�nhm�W�E�����b��O5o�����u-fEփL9�� �ֈ�n\�oc�qSH�]��E��'�}Ş/X�l�*�4��Ѓ�s�J}��o�!�z=@n3�Am������mZ�j<F��	&aj�T�����B,�-������v�~�`�.����gp�E�/	�z^;����m�bP:i}�u�����CO�䐜����6�o)(]O�fV5@�-ѫx�a���4 |��q,�_vJ�X���۔�?Ǌ��&f5H�#P������\�����8f���2 ��䐯/ +���� �v���Yr���/H���lBĞ����P�Z�$�I��9ֺЇ���Q��  2���<�+g ��Z��P��+"�"��s������xoZ�·�Df�+�rh�G���j��!��s\��A�S�D���.�[�V��2�A��J�s��InA�U�Fc�:G g��}�Z"L�B��C�T���H�}��B�P��+t��^�2��Y�|:켱��#�SYMۄ�o�UP�?�L�)�x�a{d ;o��z<{�d��������v��K�I�߇iQ_<}��Qǃ�0E	��7�Ai�zةLەb��nr���A�ϋg��Ҽ�(M�����"��^ɮ}���ٸ9�VK��:�¿&"�c�l�x�b���U�2�	Ya�P�X����d]�Zy��abE�7�cr6�Qo~��y�7V~�qogLx�}�e���e���@GQVmV�ә$��;��7�5ڴv����G�\�ΒB��_q�X�!�L���A����p���c0ۅ8-H�@`Ǻ7�G�bo^r0��K+f�N<��������4�h�^(��`�� O���RP�6ŶN0�h��p�c��A����v"�xc��ߐ�(�3��8
���G.���M�T�V�Ha~��z�����[�/�4��C�rk�k�7d�K0N��l&ً.E��OT����S8Ɇ��D�BtCi�H��7*��j�Q�G�~y�G"�o�����MY�I4[�)��q�נŝ:<�t��`X���x��t<�ici�o%�ˍ��/l��S����V��ǽ��o�h��Ǵ�k��[�������P�a _��$T���1)՘�0��'bK2�.P�˷�I�(ץ�S
?v������b'Z���8 �J	=���h_��"�q���T�0���vib�8�!]�H�IP>������&�WHV�*�[gD0�〕;$���vV�{hq�㮰�j��	�3�����A���J˚=կ�Nʮ���^�=��{�W|߰Q�$�-N���/�uGѱx�Ǫ������nu�W��	@b��y�i���L� B��G<���:^�R'�x	vc�]3�����9h@�lm��e��MP��EE:	��r�m����g�k͔k,[��`�0�!N�d�	;�X�NU���}a���?HD�Ob��!Q�O�E�t�|@�n��,���I�g{�l�NP�3|���MV�a҇� �*<��o���dLQf�R!4��.|��v�('f�aԏ����q�Q�Avb����5����s�.w�6������B��N��M�K$J�>�6� P��Qy��/��l=N�^9Fe �'̿�$�ݞ,���aK��G%��Z�;z��&�NM�M��[�֚�ߘ_h�|�|��F�,m���6d1M���,�z�W�X���o�lz��p��ᒽ�@Ϝo�H_�b�\����ᆍ|
[��z��w�q5~9N�fw
��R�����JP\���)&*���y���c��A`�V1F/՜R)����>�F�cT�jK��K?Gr��:��SbU'�[��џ%S��T�Zḥ7a�l��9 Dx�{��,<�4�
�K`Q��2�0��K&#S+g�oWS�S�2�Ru<��ʰE�۝C�=�@��"9�) c8 [�r /#b�^C�rbmYX^��DQ���/�m�N;�e	x�쫊$��}X@
�t�)�:Z\C=4�!���`�U���p:��ب2vq�>��"�w���g9l�[~�-$!�߻��>��y�v�U\�7�S��V[��&�#�A�"�cD�q�zM�fA��D��|���e
j�nb���k�Tt�9����ru��{"x�?�+�$�:��3
w�
���L�2�E�*���?�N/#���4�q�Lޔ�N:�yō��q.&�'�>#>Yi�W� y�[��/���O'�P����a�w��Z����u�LK�n�6���x��@�+��W���XE�L��R��5yq��YX�S��`#�jg�I����1���-��[7���F�
�ҥ���jQ��g(l<���)#k]kYX�ȣxE0ʚ���DM{:6�=DmU�[7���\���'VN�xaˮ��i 6a��:�C���0�`������sCN���#�|*�t�籐�W:+��@D����ei�����q������z��X1�غ��K*^E���mY;|-����K�����`K�ُ@ւ�BSɸ�}t�27��:ۃ�NS��m��!E�6��n�V��3.N���c�s��V���u{���^y��@K21&�W��،j����I�,��n�?%�nG�E�ũ\�U��i���ĤV�����ϔ�:&���}^��/�z�)�҉=�U��o�H�i�l|F��+Mڹ���N~ڝ�t���_ )q�EZ����Pu�e��F����קyY��!M���7/�U������wb��r��S��M�#YŖ&9b�Tt�V�-~�6J	t�f�U&+�9q�!�nWW\�~���E���@[�m���Y|Z�j=X�w���� ����e�WK�mĊ�l5]Zz1딄�/�����P:l`�~�<�{/l�9��k�J��K*=���_gU�ߣ��"�?�5��1�e�w^yl�e�B�q��N�86�]�/ 
aڽ�Ij��=��je(~b{]��m��M�+����F�CcL��їw/Xj1�[��(�v!��9�蜖HPK�1���*y%�uf�:����|6�_���!��ط��]����g�9�V�)>�2^ITo<�����F4����p\o%�Ϻ�μ�`������q#���3H,J�d�|fvnɌ�p���5��XT�诅-�J�'kM�^�N�c��Ň�K5�׿_c4ς󣼫�
#��vQ�b�}�����ղ���T��o70����jɐahB�Ğ�.q�븞�;f|���HM��2H�?Z����6���G�802��4�k��:���u!�r�������:���\'���l Plk����3Ak�A��$ハ�#�s����;S��!]�t��3�g}pv�	�鏞a��Q�8Q� d��Ε��t��y6������>�#����P&�L��_��E?0�ޓ⌦hP�(�ٺ��91�,y��G�Z7VZ���Y��3u���m�9EI)_S�)Yw�c�*̟�n�����	��K! 	�2�N=��'M�lۅEN@�;����uJ�:����`I�=lr�	s�. j���r�ęIY��F[?��L5��� X��\b	_;�tg�!y+Ԫ�a˄W;seq��r{�-䦗D�,�����-J�k�y9Ҹ5��ٺ��b$� �9���y�#-	h�b�*$4Lɠ��\��D��Olg�^��|�4��.}�/��9nE*6m'���|�(+Xl�v@�}dT�����40W��ોʳj��愗�A;�^P�8F��;"���f�C�8?� �)�f���5�J~�G2������I���ȑ��6�RTo@o������� �י�GX�W81��h`nB��������+*��������H��z�四O�[�=��q�7;g�������Q�!��pGiwoBy���3�Q��GOzfc�x�0����͡��Iu�B������r��:|S�z���#D��m� �%]�l�� !�b���	JHM����/t�����dDp\��젭n��d���[�%�N�oy���H:���	�Ł�m�o��,i/�E�r�#�,��=��K(7����A^�M$�:*��Y?��������;K*�Uj!�_�~���5�&:��>�tj�j�R�^4�k��Mր	1���?��<�즈���d�8�7�������W+�Ɣ�	�-��{�gQ,�����*�뽐��08�>�!r�ضZ�Y;�� ]?�/��������d�T48d��V坊m"��y�X��Y��<��w�}n�/��Ԙ��2�����MZ�V�mO<Y(������7(Y	`�a*k��MA��p&�:HH�I�X�]��1@i
j�#i��`O��*O��E;p�w�6`.&��[��f�$2M��x�{t���|�r)lK�4^��P��l��&��Y��m��A��ݠUZH�|8�y<�^a�p�2f�Z�/��U��ɷS������fK��r2�j��s1��L10�׉_Y����û�&x;n�t�/�=�W����\XN��L�R�}��l[ݼ��k<�!"^��d[��?dt{5�QO�����Zr.R����L�H���_UR%Uq2�\�xb#|�o8�l����~f*g�P������ �nT��&>��ϴn*�$����		I;�vil�4�f8\1�q�X*x2A	�W�k����^���c�����r}7L6J�Jׯ[k�+*��{��Ɇ�����g��:���3tQ�$3�<�z� Ͷ%�®'�KG;�����&�W��!����F�7"�����U1ِ	i@�2?����w�;ڲ���Eq��2��9C���at{�ѓ�����}kr���QA>�p��a�$k�̶0yE�i�'�w�g��w����n����l�"�[94h�x�.���~/�q��v���y"�E��U�a�ZG̬��F���%I���
�ʣ�>8ۄ���z��R��Q�_$�����h+&�z׵H{��x�,��&�:<����U���o����G+X�hA�$���=y�xeL��5G��5�b�����|S�p�x�H�9W��ua����E�G�����,2�ּ�Wg�%D�Sc��)��A��a���++��U�9��#U͉��X���GP�a�Z����b�r;�7�}��/��i�P�B�m������Û'b�^��|�3�5�S����<�4|���NӪ�7��#���2���T�g���ޙ j�"S�dTF~UrIJ�ZD��'N��b���!��3G7᫻ Э�>�0)[
���)��s�����ъ)�r/�8A0KM�جt>Qmk=�(�i��Y�]{�������y���G)��3�2O�fc�"`QLis��գ>�W��mn��7~��Q�J;K��z� &,�h�yXfme�xڣ�j!��5J�ߥ�{���0q�tv��f�Cۉb�5��J��1o@J������)?��C⫣��"�r��,�j��(/-���YX6gPtHv�5 ��a>��S4�9v���?�&�!dԊ�B-v�$��wL�[L��o�ہU(��:��5ϟz� �����sƚ�����K|zj;� Xݜ<8����`]��LO?B���Ԥ�E��/�x1غ2��No6�{��Ȟ��6c�I�������5�yƻ�>\�$` ����h�Of�U�&��p��-a��ˁuX��^���ܺ/Ke�\��R�
���*5��d����D����[�%1&���{�9�~��|K1x�,��%V9�u��R�lo�吂��_��o'"�����PF[I[��TO���� {�	��K~�6�M���a->�\����"pH�)���<�=���'e�Ep��hȊ��3���)_W�ͦ�̄<8�ۜi �TG=�j��]V٦�͋�i���hP�[k;%�}�Ο�������Mpǚ���LG2w�����-Ϩ�7*{�;�Y�O��ǳ�P�vqg��̊���S6c�zd�T�`�v5��i+3~O��������ۻD�I��8���g����v��?�-���48t9:*���YC�I�!y�E���F��.U���sxsy]��9�*_����4]6h�ԹU�0EA#�c�p�V"�	��bf%���Q��&#+�~h� ����ymMs�0��D|K|#�!�sL�Uy��G��/K3����*y�+����X> �x�_~8
����b*�]	]M���3I���fD^ `���j�e���0]-�}�U!7���^'��_ʹ����/�-��<t�/s�qN�,r[I@������fqI�Y|"���[�·e��ׅ�F����_�3l�t��<b���Y:���1���H�x4�;�S��g�XO�����HgPU	'��e����f?���}��4�KP>�ʎ�w�<ӑb�klБ8���.�6ścJ!	��K�`"L��Ch��X%	�-)��\�&�����K�pڜ6�®�ף#�E{�7 :.�_i����)�[}�GQ�_4�x�n��MPh�̥�K��pQ`_�R݈�K�����X��f�pę�Y0�:zX�޷[7[�U��6�����ΎV��A#3`��MC��h�B�eCd��V2*/�>�F�4or���m�ws��\.�_	�ΞcD]]��!虩S<�0���!eH6���%1�w!s��
�n�%��#�v7!�+��{J�l����+�s�X���TA(WC&x�p��r�[�k1,�5�����u���W�7��b���0~�����ͦ&��)������(g�`$	{R�;o�@t�#VEB)������i��
����H���t���,��Z@��.Ҿ��I�9�	�6���ݒ�P�F�3,�0|J�kļ6m��s��+�b�5�%��G>s�ɑ��d�r�K�d�I�G�'�.&���$��T�#_'�,�[崉л�j�)!�ώ�F��p,C��c����b��2:�!�&N���V&�S� X��Ѯ�=i�����p[?�X0��$G���;qY���B�:�:t��)ht�Q��8�h��3Q�e����ړі�&�6%8?��AL^_�!K]Y*��_�"0��C�w������
QR�;(�k�5��6���:����^v8��5Uљ�&�D�a�\T*��ޝ&�D*"�U=�ߩOd�J4��D�_�z��qGv����W#"�O*��3�t#�+a�of������,7�����ʍWKԻ�}�xF�;�F=z� ��a+Y�q$.�Hd~��t���-� �:��Y,Qk�"��t���U�I8o��}茶��YE���L�-�H����z�$���[�7��Kn�0�m^)��Um�C�W�����1�5���7���21D��d��*s�(\w��+$�H��I�i_��5�w�J�ӄ3x ���/wR�ν���M����K3!�����_8 ק⥟!�Ы�B:pG�iE�b~����ߢ�5:\�l���i���zE��`y��.Ap�VHY���L E{�1?ׅC�%��9U��q�jS��O�w�:�
�4���4!8^�ްn��3���bE�"~�~���b��3&��������3FU��A�0�&n����]>��FrbS��I�h��&��Du�(�W��v
�j��ԠѮ�4�5���\y>�;Zw>}�:�)L%��c�8?ۛ�DPi�����27|$�>^BH	��^�Ǹ���h��j�;S�v�ٖv�,�wpد�~G&შ��#n�w�2���DܣSǺ!� ��*�*�����nGS�1P��b��/MF��=�]���3����T���h���#ҕ���	���#|`Bse���.;�,�{kRǩ����l�IY��+|
�����R�ǯ����x����K�H\�N�G%e݉?A�Y}�Q��ƾ�(+�[[�*��a�ͳ�x�K���{����b&{�+��-ϕ�B5�qv����t���r�L^m�!�x�S��������e��iy�C��@�3ڐ���L�����|9�>��ʱ��[���$��[/��:wcvw���XGWѲ^{ !^������&n���rS�L�w�l�vWz��V�����Is�����*{ N����P��r)]P�O6���cr����DK*x �ڪ����Z��q��M>Wg�����&��0X�#�_����Y`|a�	^Ӈ���OS���t�#�C�4CҹK�/��`t�v�j)¦���:o�ٽ����N=X΁tQ��A�4a��`����d�4��:�g�*7���%�\1Ӭ ��u+=�B�ʂ����������C��xq���K�R|�@���j�uEXu��@+?��v�%͕v��;�O̊��99�B�{<�a�Q�>��^��ɚ?��D����o��G{P�1����n�������:�V��s���z���0}��"��SX��@��#�~W����7�v����LqC�!f-)��IMz�d���P�+�5*O�h*������N�C|VO��x�n�sԣ��������|Mhs?�)����^=��h
T$ � dF'���&�[��BJ4焘�9�>�n�gS�hh�Fӻ����|�	��D)���ŵ��:s���>C��n��x���eJ�{�k�� [�}I�auT�ׂ�|�|���] ~�k���Zo�f@tYO�uR����ia�諆F�ڌ��L7&[�VKU��b\�}q���(aS���$�5H��uW�sʪL3�0�w���ݖ
��!A���Wc� i��n
0� �mVf�*8���޴(]h`ݛ�|{��aӳ�M�3�Ԙz���m���@�s2���2���z�zqpcZ���y5R֛�l|:���-7�]��Q
TP/���番$�J�I���|�WH�z��q�����i��t���I��ӂWN{;���%�OJ��y��<�E7�(a,�8L&��1�����Z�|��GD����>em���w�.�"h���w%����z�Պ�^��S�y1�Ųy�͢k!���!�n��#�y	<��&Q1Р��A5t��|C���#�;|&(��`�0J����u�k��ƞ� u�FP���$#��~Z7z����ޙ�y6��9�$��;+�v,*`���1X�r�!�4ckR�w2k�?Z��1���$����<'�n5(����Nb�
c׈����s���F����(g�"�k�א����n����h?��^2�1�4J�H��l�,��fkĄ�5�;S�4���M:��If��έ�5~���V.oޜ�@�6!j�G���8������m����~cM���();�}<����m����\�G�}�I���j؜����>�dn57r�8����-�b�������l�Et|�V�q����kv ��m��P2��P`��:�J�����ϡ���5���U1��|��z���T��e��_&�aDJfNX{M����W�Wn}u}j�-ģ�uH�Q~���,����dH��6�g7�T�Z+��X-��x����f:z�/�@ʉ��f���P�::7֖��ۂ~����V6�SRޏ�ce��ӌ[�
�βg��k�|�㌦�����s�>8p���5(�ӂ�����B�I�o0���,s��a�xU	{���!�H�8�N���V�$�'���M
VO�ˌ-)��	Q�-��p��Ļ���)��ɒ^|�
�
8��G���	9؏�w~넱��K7��r9c-D�ȶ;�W~s�&����w�¸��J0Z=ӑ/���	���e��v�`,gO|�1b�4�~�*w�7`��V� 9�tx::x�g�C<���&i�'~��,�9���MM�f9A�DL��9�g�e�b�R�	���J5w�W�h �>�On����D�k�B�_�V�٭��t�ˏ��z�I��A�K����y����PK�Te��`,V�)p%����
ch�+sQ��?�}.x���Y�(���t i��>p���/��1cT���zv^�����{��"�>��%�:�s�"�B�lBr�Kt�A����l��?!F'I�"�bŤw���#���,�S�"YK��s��\Ŧ�!�����k���<������h]��ڸ��u���9fJIMk� n*k\hh9D�4A��؂j�����rB���{ k/���g�4�@�a��V�Q){bșe�D��_���������;⚨���ܾd:��S�ř��G��N�d��9��X�7��� �ol�3�R5���,����m�ij-ő�F�ϱ��b�yH���<k�u�/� p���]0I1*i2��3��C�Q��邧r��s��,����*½�41��mVs���Va�ۘȰ#�������Y�~��[,����e���^��;��m�ɐ�d[V�?��fO8��s�֓�'�
����FB�� �rǭ�gYh��a�yD����q~���y�*SAR�f�!����H�-�+��"���%�ZV%��M��8JrӬ��v_Z��$�\�Ude������Ě��R��g#�P�f����>�G�nN٢Z�}W�	����t�o�x%������ڰ��PW���^�}ڌo*� �`D�mV��O���Uy~gP��_��N��Y�(%�� ��vY����ꅗF>q
���R(��m��t#Q>� k������V��@)HZ��@�1��n�F8~Ď$���W�O�/܇w<Ϧ�r"��2��L@ub�'�M�\����7G��'��̒�9���*@$�f������31��7=���� ҈G�<�П�p�.p?����Q�>hU[A:e��$L��om�u��GK놴�08��R ������0�s��2$�1�Ɩ�s%�dpmS/ӼO5ƾ�lm���z���N~sz���a8�d�{�n��h�g~��2����Zd���@�v���hȲ<�Vg�(;���˱��7�p,
N\.���?��L���S+3��&��~��5�<v2}Ӏ��.�0�_E�d�&�����$Z�ñ��|C�8d�:�u���u3b2w�V�#�c5^�����	vrj(�~T& �Ȗ%;�f�w~oW���F��ŏ#2�:v�un-bF�%�\;������q�;���@#a28�<�<���;sZ��r8:��F"���D&<�F5�T���M.IC}mzz�w�E��b���m�4��.�����#��Y�1�G�SR��*��t ���*Q�bx���Zk��& �&`S�x����*EZ�����!�k�7��_���Gw�_��Rk��|fa��E�0�ߎtF ��ˈJ=�?�?�Z
l��������(�.�Y�^����c'��R0&o~�i;}Ѐ�vQt�WI���j�QB��ݒ�iɅ�9t8r�f'�����+��>�!G��{�宧9�s$��Sn�e��<����U��������;0�7D����a�[2�X�^U��c!{�q
"��h8V�N�C�}���ۙ�����|˥���^�c�9���5�3ߙW!��X3g���D���@����3'��K��V��_~�p���Yb���p]�:��&¬�|������X�0��<���y�����l�\<FpG[Qp��m$���H�7�A��&Rh�q�*i106���?�1����>�-֙1��t�'[�)��^خ6*a�Y�k�S	��e�^և ��E�zM��ssM��D��*������O:Ԥm,���ZF23�z�5af'ϗGu���6}��ϲz�;P@ q�j8$"�h��ׇ�P�K��RDu���N��+L��mҸrJ�����xvQǐYd���H�p�e"�+�q�6�۟>ns�͙�W�[��=v:7e�2�rX�~GD�Ŋou����N���1J7��Ã;��|�oR���{���ܤ�V�1(�Ê"��1 �I"^��ZFB��[Ѵ��m�n�x�����3/���g+�V��~j����V_2 =�ׄ�͢� ��ZC�i8@�"��Z�0��>�ʗ.��]3R��_���?�At�G�����<�J�e�n�7k�'�	4�'FȟG��5��B�`���2��&�};c�{�����+=��v&z�����~]nB88�������ݣ>i���ú�_�_<c ���:~4�?a���m.�Vc�ˮ���� 1WeN�RBƔ�J'>~d���=K e1��� d��ԗ�Ťt%@�j)��`��ӗ�ǳV��f:�igP �����$��=1����~��r�6�E��P��ʾ�4����e��u8K�u$j���@����x)!%���-�.I��8x�: l�u!�u�2Ϛ�8N�$G�m�f��u�c�0g�M�>�����72�O��5y|���A�x���n�~�x�Jݻ����g�DB9H�ܟBid�b��*�س�����z3@F�4�熬���@2PL�����sN�7���ƌěֳ���5����]젢�+���e�'���<�y���$�z|yc�I.p2����N���/z}CnR��U��nOU�)�9<��ح��K�'B�� I�AU��w�b�U�]Q�)�+�r�f�W�]^ ����Lt
`��&��#�{L�����j����K� ��s���c�M=��=C=pތ�5�r�N�?���w�%�?9�h?���J��E��i�#C$�빈l>�{!/a݉xFM��ik��l����@�����~�
�= �����������4�Ư����eK��~'��)���K�jQ	ع��N�?x�X��-����6����h:�����=]C���l%7�-�k����?^�w�S��;�7]$i{��U��yB�|j�����>8@�)ղ�f7/:�Iǖ�Sз�9��Q���ᛰSe��YnZ�]f��9��r�I��HH/��M);]��.�w������!r�b�b���iB��:ȓ#���,2�[�]epdyMfR\
e3��߽f�h�x��3*;�
.qRC��I3MK[5"�_䅘�s��o�Ii���M3G�H�q�ݎ�e3 Ns����>b6M��~{U�8��t�C�f-y�nŠŒE��c���~|�w�ӟQ|'n��Vuo���H�4������O@膌E�IY�]K���-Kd�}��gA��+�I�ʑ���Md����U�qz/�o� @�Sw-#��'
ҲZ��;_J�.p��)��梅�n(�z�):��|�!$���a蓲mt��q���=�m�����U
+w��>� ��gR�w�j�\���}v��L��H^�Qde��͝Z�&C��uI�B��܇�� A����� ��	�����5i���A8M9��0���X5�d�Ϝ�%���hgk�1{�Q�u�L�?�:'�6��#�#{�}
	-����;/mB����*��?��_���(^�Q����+T�BN�|6���|�S���B,oD��Lґ/�-*��X�q���h��dy�Ҿ�G�������!҅mc�{USě��M�x�y<Ul�k{��tN/�j =N�{��1��ϙa����KG}�$�SxDI�;˸L�{̌^`֒Ysh�Z���d�g2U�����߿��yڟ/b%��~�[I̩�EB�[����Cpy�,�&��-�n-�+�ꭠfB��^�߳;�9;o�g���tW`�}C����H�T�|�7���&f�heÅ�ߺ��j�ep`�(����(��������sm��U��y.ʢTO�7?د�¨��N���;�c8�`�p��}��?�M~@���u�rl�Ӷ��A��V>é�^��N����S�~§�}A(� =(tW,����.�i��1��,~Nu�"���c!ݵ,���KUo�����ܬBz����C{�'&U2֣�x~��͢��վĊ@�IB���yee�] 	O���b7�A��O��Ѻ�3m��M�������}ŀxY��&/�?M_�o���:�7��%�H��M����S
�b.�%� pQ�ѵ�?�ߛ:���lRLK�IEgFQ��>�о�p�6�l>�$f,k�z���inğ�H]������v^=�ơF��&��h�R����WC����jMX�Uv�X���l}�Ɗ�YS/��1{�Z_s'l�B��f7��X�(xuY�1��V���2�L��Y�P����ig�l�%��-��C$�/�;a��)i�M�z���Yש�,v.�j���̗�C�y͛q�ftމ�Lq-I��	����n,�@2��ӳ���$��]�hV_4������h�:(�e�@��n�0������S:\[�3C����ݩ�7���a;um���֗�&�ڪJ��j���O�ty37��|F8]ks������-;mh�D��:�+`qQ@�,4XpǙ��*r����0z�zk0�-B 3������4��GSQ�_Q%�+��oV	�/J�=���7�__�T|Hk�2xf���a��:�nT�a�7�{���@vaDG?ە)�_S�1;FU3m���m)�{�]��%��Jӊ��uUP�%����?}����g��׫��9K(�`u)gʘB9�&"3'��q1>-��̛�\y�\�.]#0�ʹ>�e���W�y�j6�sgX9�>�YCPK�(H0b�_]WbF�*� J��	rF��q<t/I�Cw���<�DB�쮏�$g��*�4��9�b���!��,��`���[KF+o}x�x9�2:00�����\l"�LL4M1�L5���wS:]���e=^���^�ޓʳEG{�X(�����Պ���On���h���{��{a�W�d����i t�{���]���N��6�U�kQ�*y��9l��7^~�?��}"?�c�W�� xԳ �X~c�9�L��6���}����n����H�a�|���F���_J@���`>��ko�V��m�]�k�%��O�?�)���Yp��NTq����D�^A{YGq� B��B�	R������I÷��ڡ~KЦ�	U��t���Y)g?r�����E����v�A�t���J�ƺ
~�~#�ƙx��U�,j�s|d���KG�7#d����-HkN��g����50�.�@���flF�[7����%�G���K[�L"�!�L�:�qS�Vr_4w��;���e[���
��:˛��	am����V� ��S�9+J4JLg����HrXM8h��{3�K�@T�FԚ�~�>O��a��{.�r��bȬ	����s�R�3�
�Pȸ��յ"sk*	azg^#5؝��U¤�jEZ^�/���
@LXC���& ���I| -l���im� �F[,���䚹;�N<�AL6Ʃ�cjy����-: �7I�I��T!2~Mku���/�1�Ϭ�L���M~�^��	�4av����Iƫ��| ��b�������M���:� ��C+�;�Et��u1"�Yu����^��j(��n��Ph{�@���+\��A�����:.m�� O+L�W�;���������5���ǡ��	L�ߓ$b��k��m���Sn�� �F). �`~��l��y����@mu0%��X%ꬲ(%Qݎ��?9����xmO��H/����ѓZE�Z%Tmr��Y�^��;F���a�%;�,�z]�{XQ�1޿\r���@�{"�hK�C�b=Q #�k/��3I�4�5&��b���©�c4�NǢרxpfםܙ�2�@�a�X�C �ugi٧���T���̈AѨ�;�iq�	��)�)����m��{h��.���"��u_̈���q�� ��h~U�3��u\Aa�-@���G���C�8IY��V��p����ѯ�U�.m5���,U���"g"�����G��n��^�����~�F���9/~�mQ�8���0F8k6<8QI�O�����B��$�옒��L�=6���ܯ�eÓ�ǁ:�zc`:dH����A8'q�ܦ��0��~gN���Q�k{yr@��*��|���l}~쵅	���R��ZP���Oޢ�`�D�{�HQ���ƈxFX�rHfn>�� �tlLj}n��\f�N/��9Li0d+.�9�̀�������?nY��g�n�1Z[����g��*2�#�����R�7�)M��.o����Af�]��$�����GꝄO�A0��_O�vO6��a��D��P[��q��s��t�:�N��H�yR�U��75�� �	̇��(R4�7�j
�7Ȩ��q�M�8dt�V���E����� ��m�\�@E@B�|�d����Ȕj�7��A����XO+����cð��l�M$�~`2&�7�����{M��g��<(Q�������+�G*⾛̧� <}p�g�c�bvb���9~��44�x�o��砸�������p��e��h��<�Jzn���(���{�U2^�;y`�6_���n�I\y6���3=.��6��M��%`�]�Sڳ��Z�������g+j,�X4��d���o8���(��H7&��^���W�//��]p|�?gV������ě�U���r��ꎭ�l�%)���go�I���6)��h���l�6��)���1ig��@��V),�*m0���qFޞg�K���5>�LgW@:����Wg��J��>�O�����.�� 'j$
��:P'�y�~� 8���kK�@�.�����I��1�K�*{�����g��B�0,��|	1:+�;dV���n����U�d�S�lԯ
�#;����j�x��
��� �2�L$VP竨}���1�+�l�R�)�`�b�Ԧ����X�u;�6).��-5+�xȸ#$V�.�d�%�=_�e2x-�8� :�����>ѯ�����kHT�J�V�R�\�cM�6�X��4^@S���2���8[�0�=%�|@ L�g���FS���ՒY�p��)
G���e&x��9+[f��M>O8����Y����jzY�b1� ji*;�ϻ��%1�A0ؠ�e��r��E��a�!�AU���Y~��<j^+
G03���q�2�v��
��Y�.a�@�.$�LC��` At�
����	{��C���zH��߀�&����L7s�S�
��<�R,����r?�Ȩ��y�#�b���Wެ�|�0���B�b���·�{3�"�R9pC�%�Z��!���%�O����1P�oq�J޼���HrK�\Ӡ�T�ӌ�r{ =x1/��v:��z�����&wFt��n9-6y��	�H1j4�}�^0��A��Q���Uq��"#5����-�P�I�G�B9��P5�s�O�v�G�^�IT�g�ڊW&+�ᦚj���	���/�iq`�qx]�@|5��-�`�2]�P���1�x��10�%��v7����BcQ�=񝂾.1��I��?oR�ٮ��\��������8����f�7ʂ��1w�������^�ihN�n~E ��@4,�U������\����a�̙:_����E����@Cŧ��J��J/$�؜����:��C�_��,����ʞٝND�o$�Ԇ"�r̷���R���l�:��s[&���e�bZ�I���+�}Sۿ��Joi'Y���Vm�C�_���Il�*��S�<{2F��ME{��q �ލ�j��P$+L�:2��G��rn�r��y[h�V��uC�Mb��A��P�a�0��=|l�Ȼi��#8�N�}��7���������e�6?A�c#R��t�*�	f'St
�Bӱ���<q�֟�������_2�aiʴz]��t�4vv�pAO��50��B�MPH|j0�������2S:˓�<x����Jat#�t��Щ2�@_�jΫ 9��a0b���1R<}3��Q��8�e1S��g��H^���F�f;�N� �ͅ�Ҳ�.'?�sf������2G����@9���E�}�{p��ĕ8ݤ�[L;�d;�Ŗ�e�sSc�9=����fQ���ȁRݷ���a�ER|�� ԋ!vQ�UM}�x�S��D�� F�t�ZU��>��gjX]�(ʓ��UR��t�	F?搏�B����=�?ݞm�;��c�F"i� é�ǲ��%wm�;�N_9�뜃��s��"�#M�6"@�Q[ʤ?��33@�80�]k��\�������<SM�����`6����r�}�D�UT�L�\�Er�R�p�G(w�?��~,6&�F���Ň��������!���/ΘsO�C,�6,6y�#��q�	��}�@"&��G��:O�o,ʙG���>�{~��g�ś-�Y�cY䑵��l����/�/ArK�~­�����E]8�s&ZՐXi�?�:��i9p[�e�{��]��9�d�M�;��ј�jh:P�oyMT��.4&��#��P�O�>�ǭl�X���\d d� �_�Gau_[��5�%����λ'����O����������g�$?aw֊n �:����S��3I�~tF�����<�ɱ5UXɢWliV\-����K�C
���6��>������~w���[�K��̨������b��!������jd4յ��pwS����>��e$��ʔ��I�3sv ����d��ghZ�ϫ�_�F�sY�J�S��~&+�mVQu;�G�[��Ŕ'6R֑�|������$��FM�>�a�w�*X�����c`@,��aD�o���}����.�Z�r'%�T
}t���	4�4TaCe����Cu�Df��T���Ƀ�1ã8�$f�o]>:ա,�3^�q�+Z��Dˁ�� �*���'�[�u��{3�Dxf_�&���������1{L�V�"�6� ��:�3��S�]dc�d
���|��ϰ�w�q�S ��Ջ�T�x��� /���b��[HS=9�,�t
d��<���sѡ��z���4�'�g�K�S�S(lx��9�Ƞg@0[��j�T�p ���3u*�qӖ�~�d~���2 M�n�v��9�D�]N{�'x!���+97>�"�BR`�A_�^e�~��M��-:�G�[���|6?�l�p������%"��{2��i*����r�H����h��~nu�*��v�m��Їi�Y�mq����Tt�׈�0P�;�[�[��;���}I +f��Â�a��c��47�BW���^!B5HS��tT|v4`���L�~��ӏNvw�z}f��~�δ)����~�C-~Ȗ�?,Ү�,] �آ~�����|6�e�O�H��OZp�`V^J�5� H���[��L��Zt�x;�POK)�I��l=��-��(8�䪒#Y������v鰙� ����9]���?�H�i}����d )��8����v�ea�KS�dK�$�@c.�ߴfqǱ~6�q�<#mb������V��NX���)�{r~�>&�)�����_S�^��O�r&?;%`E��v�����fk�����gzp�K��ݱnT��F��!X����i8(�����������}��'�Rf-�JZ�(�Y����fձ�3��.�jt6�����g) �m�OP�`�NiH'��������g@x�5؛�r�\��l�'q�H��^:�l�'��9QU1���o��4(6�uU9��+ ���2�9�u�i��H)%wE C#���:�L���,]O��rP$�QN���`v���2U�3z�=b-��9��U��Ҵ��.�G��txgz����V�MA���<�XQA��N�t����1�,	$#N�� Ӏ?2�rR��AH�V O�uB4K�(��g���a�-��S���ǫi`��<�HS��g%��d���۳G�Jz�XQbUR����I�V�%����r��C/yOV2��&�%B��h�k����g���;�fb#܋ŒOW��S�5�p¹z�E�}4T�u�4�Xk��[�-�H?T���KR�"∑.N�$Rƫ�d�t��3�3ƿ�޽-���s�rKװ�(\���1i�wҍ��
)�w��(i���f,��9h[��eA=��4���?S��KrA��E��T��'aZ3���V�\�>!��&��8;|Ę��.�|�%EʚN��W�fQ��уG%��AIߢ ��)hƁ"�p����RuW�n�-ß���H����3��n�kc�Cf�V�{`�o�ck;*^gE+�:[W�k��ff��K}���4�E����r[/��ӆ�Y��`�&��+�&�gM_�l'wFB�EE䥬�,��I��nI��vEA�Lϔ����='����RRg2�q%����m�e���_n5�/��S�0���
�z��d�x_�v���`�0׮�6��M����C�|зy�}���I��Ĕ}�=��B��:�Q���0̎C�,jM��ՙx���5P� `�V�M�F�>!�ЅQ\�O��/nN�� Ũ�������5#�\�4ѥ��%��&��<���+���L_��j�;�C)}Ӝ?�͜IiE�C6)uYi��NW[
�x�^�~�P��KF�����;�Dօ
�B����C�ԿY�J���EV~U&�znS)��š~K Q,�e�i�	��~"�ք��ȅ����դ얂P-��"��a�	7�J@���"�R��!�#7�F�2��A�neXΖE���K�%g� r�t�	���礪�+�@`�B�a�nl����U�f(-��s=}tX�z(�u �4r�Lⴌ���~*�Z��lU��]g5���ܫ�zȬF־��g�d�ƬB�/d��Z���^Y�S'��Ͼ�K��31�R�dЍ�(\�I>���1Ә�Kj���z�j5�F�Ԙ�:L������E�x��@�\2rɕ1�x���s����d4o�Cڲ��5S�f ����GWPI=ܥ[O���7��*�����Lor�5
l��H��O��&0x��G�:�d�g0mEe�nW�.�>d�Xht����+| ��\]H7>j�3vK�i�1g�X�6NM6���Sp�q�ic"��,�i��	6>qQ]ڛ?��q��:=��J]�������{F~K�z>���4J@�CP���[�v�2�1$�TAnT���k�Z�c3����s�*��~�����U�i�F��/�t�+��4�(��uz�j�r�c�g���������k(O�;s��q�>�t(�$9[󽬜��ƄB�u�rJ�]�xF��3L;X��%�K�������SP�����b!��%�g�ؗ�/lm�w��^Wfx/c��3�KQ_�HPvVv�\��5����<¤Ewp�}�pX5�?`��qc��<�$k�) �&�_a�pv�X��iG�̚��� 7�h5�d�:�{��\�:�icH�z���h�\�M���&ͨb.o �C&/(O����M��,��,��::A�Ҕۙ��i�&A���Ɇ��Ń�n��AX߁ ���+C�]�c0�4���N���H��%}40V���
+�}vf���O�0����x2%��bFN�.�7f�X;0m$����A�,���Ɨ�Q1;Ϭ�����`9 y���.�	k�'�����i հD~ �`�Β��f��o:��k�*aǌ]���џ����k:7�	���;(丞�<֏�ޠ�g�Ԅ�y����DT�xH��m�l�{B�ӌ��c�݇��F���j|����)���6�@ ��;��*�C ��J�y��5K�AP��y*JQ��"����o��Mu�)���s�aiZ�	�Z-H�3Aj�[E�o�)W���$H[������=��,�rr�����szD~ٹ@�M�g,M�\����$�p�d�g�a��hDBx��X5�GR�X��w�����87�>j�g�'��Ѣ �^�4Y4�Ľ��kK�;�YR PY��bc�3�ê�e�6��_��E���uEX�i&�yE�39y`e��v��0Ŭ:/;89[UD�Ґ�X˨Y�s�:C?�)�C>q}PW���AΩ�ܒ1頼��N�-?Ǜ�@q��0vP�����O�6��T��l�������H��iTCڷ��+��v��q_��8E	�OJ�:�Z����^2��"��fB��CΎw�RR-07t����@�J9�,U$�g7b��kL\6Xدg�t]�S*g�Ë�����f8%�4���#��?��sP?i�+�5��q�t!��0wP�+M5T1!�ǟ����?�gpEŅ�vw�)=j�X��MA]]1��YB��^� 
�
������n`� ��NX�&�+�a�5���v�݁〻�>w��3b�� �-[Ô��<��g�3p����ߖ�A�m�N�%;�sD|�@u��*�W ���������U;-���2
�h�A����Ma)f����my�>�u��}�1t(��`��֘�˭�}"�v��ូ�����k�\�	{�>Ӏu�A]����Z����v�	�>hIk=�H�t=$�p?�p�!S;vg�̙\�u��q.�g�T�
g��E�(�x�b5	aG��S9k\!y=�3k�X�N��c\�F�+��fs�{�Qc�?n�T5�d{��,�m{���bL�+ϫ��к��V��x�_�_n�M������3�B��>���*F�ZA���$���{����F�ބ�h�\v�V� ��{�Pr�?u,��N8&�P;C�ː|ۥ����c�ތ�Q��{ݹp����� 8��׊��z�����mEٙv��K��s���:y˾�����dH�|��S���/~�DR���;��J�	��n�7
a��������/V���'.�w0v����Ld�(f��=Ԛ��[;�gһn�U|��q/@	F_'$�Q�Ȯ.Yf�!�V)I\�4�Г�V~_�!#�|���`��F����s�Q`�pMջ-��F{�/�B��Q=�����E�?�'D�'OƜ��W�x��{�~P]��Jr8&���ް�`P�Ƙh㽺s�W��eW`�C����
td��̬�_;�e׺�d�Pc���13��r�Ζ�-�u��N���Վ=a�K7K��\RAl��΍$u��R]G;�^]��M"�7
N��o����
�������^�I� �tu�J'�:@!�!r~~�2&C�2�P��C��(���ʤ��KOp�V��K�`��ź�pG�0�Ec���w���Y�U�ء��`�[2��F!��7"�M���&r�V��![<��3�f�ͦ�Ij9�hD�uV v)��0�Lް�| �h�ugrD�JO��P_(���4r�ܸJ�4P{z�@�W� aj�t�O��2՟�8���²N���y�e����+��-��CP��(7Ɲk/��Zީ��5"iQ��u������v��z�-�o��aZ�W�zh�L�	�f���0Z�LO2B�B�7B�E�x��[�d�[�AW}�Vd�f�0K4���^U ����PS��	�Ί5'y�����/�0�Kkr�1�>���7�h�NUT�z�K���r�(��3v�()FԻ��$��X���o���ދsܧz������t�IW
�@ PS��Q>�k�H�%m��3�](�6�Lh�5��l$H�$E7a�m�^��7?G�����YC��x����A�����H9&���c��)�"������~3W�*�Z6T�ٞ�ǔ��Iۓ��5�f�5}m >�@��-�d��@3����|��b�E��̦V��Vv[��x>V�H��=�u�v;�����A8������~�9��G�#�"����xp���@s_ȧ�@�~DJg��O�Ɠ#�\��p�c+�������w��MgE��t��ç�����t�&������t�G�$������~[sy�� ���VE���9����L���T���*V�d(z"���\dz�E���̺w5A��qzu��j����h���l���H��K������er����s�
E�_[��8�O=�u[��	*�B������sD݇�+q��R؞�uw�0��r���ݮ�fa3��v��6r�:3�:���Q��̇<NiѠ1��}TSM%�E�g��"��{r�(�=��A
Ɵj.|����fv=���t���T�
TN��M����Ǫ����������a5˕!���=�t��D�XY�!�����R��	����2s����Y��@��`y 5YEݏ�լoh���`�
�3��[)�cmjR	�s0�*��[L�4�p4�M��ˀCR#vЇ�`%ia�w������Q�M �p)������Dh����E�ݱ@��KS)��R���[aW��Fd-K�qd8�D���`���&����=lK��x�J��gc��T|���H��~s������gV��R �+�e\���i0%���ɮ_x��;�.?�#f�UF�Q��ǚfs";��@��=��h)jv\�(�ж�I<��۩��vH�G�ޯz�` �ގ���ue���=������������(�k�`� M<��2˾�XR;���)�ȟ�y�\Z%�\0��'Es������_��.˧K��� ���	K�ҡ&N=�Eh�s|{�*o@�X�������Z����Xֲ���)�����6�m��ɡ.M��2�:�go�B��:W:����&KP�C�7������O�1u��t{8���3C��ᔶ��,�W#o�߽ȁ��B\������B���YԄ|Y�@-�_��i��-�	�h���R#�u��,đ4U`�2pT����/�D'?#�����u��ӳ����i�V�e6󊛀)s_��f?��I#tl�J��=l��#���'	+`]�!����dPk��%I�t�o�}Ȣ7����Y��� mS����
�f+�B�$e͝�Š����U�WM��>R�<�i���[����=��c=�0�p`�kI��B�!���'�i�7j�=~j�;mZ��\J]������H~g��Ny`��N���+2��S��m�cǤ�i�Ա�rL��4[�unf�̛
�f�i3c��;�w��a�v
u�"�#j�z��Av�:�oSc��9��p��>bJ�	��;���䓭S��͞ST����e1�&V�4����s�y�&�ʪ���e�:_�xϸ�3�u��aN��A��vۯ�u��T� N��L$�+L���6�4�\S�{3ȋK����G�{Xgw_A<�~l�zEmE&"v�J��*H_�J$dJ��<1C�v����E�x��?���-tÉS���a���bm�$�B[4�~��=X%s
�����N�.β��
W�9�-7o]���3�D��V!�	�z�V6�������h/��v�L�@�H����Q{j����Z���o?���'uu�t��̶���N9�)}����~fשi���Sr���N��
�{n������ �|���l���vQ���y+2P���]�p#��^5Ě����Z��_����#6'n����������=�q�~u��\��R����(�
�j��T�R�r�A�]լ��#�¯����T��߰��Kʗ�w�+�n{�� ���:9�?=y����oҞ��=a��m�lp�:�>=��jUk}��.�?	Q��eB"j�!�&�Ts5�|��`�jKhÏ���5���y��۞N8Ζ�ۅ�Kx6 ���6;jT�{�_P���W�Lo<�N 4� Շ��U����!	��!R/����Ui�����aQ�h㨫����ի��*��p0�	��������l*a�'�3:E�8����w�z�ǔ�:mY˃��1҇		�ơ�
���$ۜ�x��A�'h�>��h�&�/mf=¯,k����(��A|�J�9/(s7�$�h��|��Z������)���`����$��%O��=�u]�|Df����;�B���,3�W�#��S�nK����jl���s��l�	�u��J�*o�?C�%uF��*�P����Z{a¨���c7-�B�93O|����)&�f�5]�.��Z!�Q̿~�
�j��x���Rf�T8����7��d�G�����u�,,;k؆��0���y0��~JlHeT��H���ޡK3*�K=}���$75��zw�vX��	/w�$�~O���έ������o�'�W6�jҪ�Xy�;e���F��a�u���`��8��BӳܾW}
?{�rc6V�K�����L*�I-�9K��w�������T ��d}0�T��z/�����͹f��]���� N	Jj-[�泓Z��_�?<`쎧�Y?L���u��6	s^��v,��M��1��'YK�1���}�h��Q����vK�ok��"�$��Ri)1ԶѰ	���T_L%֮����ҫ��e�W�mAgebļt�0cZ&�#�;Hλ�V�>$W<;pܶ$.��b�Ow4O^7�0���ߎ��{���D8� E�Q0������:��'�(N�:���XTKBg�%�:^�F��K����0R��s�/�<.j{�l�;�ެ�i_�
��>&��7�E^�r'�L�kd�\�zA\ �}���d�����2�Pэ'�e�ۺ�p0�7j���X8�6�B�x�9ɦ0K+��X�Ze]H5�g�(�tj�q!ID�6� '��.�cqa(y���;��+
��e�\�����L0��PG��dn''��](���X!+xTڇ���:��1���<%�Z�6��I2d�v��|�vv��&���r0�~W��7 �\,ܟ�A�K�.�-��Q�!���V+ɫBE��\���!�/�PHa�Js�d��"�����i�v�3��#߀`(TJi��2tb��RcZ��(}N��X:��l�����j���H^eC�%x}-�*`�ʂ�������a��Bh�k>P�F�(�j���U�����D�_�sp���:J<�к`��{D#'���-VbG�I~���j�.��k%�%�Q,����Q��Wnx�z�Y>dP����D���L�i^�#��u����)9CE: S�����Ɯx��������i�,�����هAL�yܪ��E��YA�if
�vG�l��l���T�@�[��s���ldF\�����'G�Y��w{�����g��������=�D�v����(�W��]u��Y����?�=3`�{/C������q*׀�,������>z ,Fl��o�@eg	�[.&����es��,mf�r-�_�Ѽ���:��g&����L�`&�)w���W8X2������F��R��Q�U��
���j�/fLI������gx&y�.���w����)��� O�7��&R���n���O!�qf�N����&E�8��
��A~1�"� ����:�n�Bac���f���"�ۜQ�Xs�]��i�	g�5��G����	M�Ҹ�&��ǫ�4Kr��jNz�Ri��IA�����n�e���V�ԓ\�WTTS z�S�7A＼�J�(oCh&V�@�
��dc�q��
Mv
{��t���P���ILU�F��tf�c�䇑��-�LMli���MG\�bf�/i�T��q~5���>��zyP�<~�_v��́����Jt���Y��"�ڵ-I��·�NP�c��5�7ViU<��Z�Z�V�1��W��"Gnr5����Ӈo~xGQJWE��O h��Ř�R��%���f@�~{MN�r2K�	@�i��J�̍�� Ԕ�CG2`z�e����em��-���(w�z���XD���|֧F�x;�TQ?�lv�0���Z�6ȳ�l������h�a�e�y��S2M�8��s���a<Vgaf��\�,��d�6�8�������a՞��5+/�x	%^����CX0x�,���k��S��d�IL[�3��Ǩ���5����Ҥ�|~����-��q���?{��>
e��-��M��
s�h��[��d ��2�DC	�c��b��Kԏ�b��u(m�4���6���K]��w�ہ���a�[4�����pL]>��^��a�h��)����x�#��#��� 1��7{�{�����(���H��M��	+@ج��{#�~�Q� }'�0J�L�D���j�˂"��z�B�Z�	��Q��3��n{8� c�l���)�#�y�L�M�9��26.�s��*܆���k�ߝ��s���䡪#�d�0�y�=����i�xmsS���r�kt���,5t#����\��tsx�HR9�|���Q�M{$����U�p)Vy��Sɮ�lIِ��um:�p��(�@-&�L�	��{k��z����>����I�v��rr�P����V"5�4"��3���{�D����B�u��R2���*.݇K�WO��N���4�Dn��%f�Cާ\��d���?R�S4�ӏ<�g��q��Dr���|��9��5A�y�q���!ӈ
Kj�5٩�e��u%�ž
����ءӦ�0�~��߀\K�\[q��C'1���qA��5�p �tM��"h���|�	B�-5V�&��m#�T!��bK��Z7�n�)����* �W�xq�B�u�`���o����]x�Z�k�z�n�ޓ�#�����D3;88Lޚ�Z�a�Ѱ��U�Չ#4�֔�Z2��6�Zġ.�(�{発�tj��Jpu�&K?I6i��΅��ZReU��$�`�z �l�����L�m�n��Ȃ�Vd�$;Eg��f,�}y��cy��l3N����1P�����3�"ZK����7gS��)�
�9�k����6������>��M�������������qC����n�����s9�7��h��ވ`�~ޔ�,۟l�(��?R��*p��I���z��n+��j�n2ڬ�u�%
�Y?��G]A|�<��F�VvŁ��ƨ����'�}kY?��`�oj�@E�r^���q�թC�(��f����CJ$IPT���o`^S���~���gz$�)�F����X4��E,�uђ�t�F~�D�E<�,�ٳ?����4�!��D������p�ᰈg}�GQ��m0�ܦ���Ԭ��֪��iBi+~j�-������#���*�B>��,P��\k�)�����v�,��Ȑ�a�c�Ҥ`Z����?��}܌ū�M��|��׼��R�gR5�U	Z�к{S�lck����I��̱�`m�؃��\�0հ(��=T h�H�����J���'���|e~��ɭq��(���K���F����?��{�)�~�^pI�K]�H=Ee��,h�b�vsk?$1B*�*�j5�&W�������;Y�⁦+T"3>�,��\}G���PF���Sb/n��G���It�A����%B����V#��%ݼyGJ?/c�^6l�p;e�y���`:�r<Ӻd��k��D�f���6�9��*�-~W�:�F3%w�!�@a�}��<v� I(��k*&�|��R��iX�"Dv��MRg�
�vQjH+��{cv�k����#���^s*�,m�߭:�]I7ܺ�^B+�,^�yr_&��ip���B&Zg��N{��H��<g��{�i��#��uRk�Vb��uZ�IS����d('�c���}LC���>���m�C�e��N[x �f}#O�R$��H\{��#]���Ɗ�=н��Vm�R�K��胰6t�������r�h��<:��x���	���I�	ހ���k�>��^�� ���Ii����xFa_5�OqD�A�c�N���3A�{�t�u4��cAeR�("�aQ���zGP����X����<	��F;���#Zє�ylN�<Hq���:��E����N�đ餷����V��"�S���d`b�,!
��$�;�Q����hh�$�\�����������oۅ]�LL���/�ˀ(c����_֝ 
X9J�ҭf�;��a��`�4�ml�\�9b���jӋ�D���aӉX��Y��\��x��,�}6��? �f�<�9�ehe�$f�x�o�5'�
�P,��j��${2��6L� �}g�x�6+�TrQ�-"�b��H�L=�J>i[h����P��^�{s���I}�U�T�I�="4]8Tӕ�?�c��q�l՛xq�c l#�:�ѻ�[S_Ķ��,�����a�l�sU���oOS)>��TNa��T��2�=-c�z��¯��ٚ�Fct�M���x��ȇm�k�V���y(5��Y�ᤃ�'rT�Ls���Wb����fR�<m>U��������eg��DY�B�C����`sQ�ּ]D����C��i���4�I�k��TN��=�� ����T���	Y�7�TD�D7�`=���#mk�D6}u|�%nm��{����
�m�N峃��IO�a�z!�ZBl����֔���&����&IG�)H�W��L�,hp'�B�����3~N����O՟�6CK�/bA�Dv
�7r�"7���4P���y�e_�kA�%�j�*b�L�յ&�`��w�@*� �S�Q7xn�f'���x��q��$��%���i�5�j���Mm� �1�*x�gK���r}�Lc��YL�<�Ҵ��?|<�-�ti�YS�.M�	���-�bi�,L����9}��Pg	G.5�79�E�jv֫�m�-�+��F��ſ֛G��1�!�H/�ic�l�Э]�ж0$f�����p��{#L�v.T��7�m�s��}ɔ8��X�i�Ն��5XL���L��r}H-¾4u5<�q��X�b��GD#��;;�Gi�"3p=޾�4�F�:M�>F=� ��
��ڵ��wy���t0��#Aȗx���g�*MEu�ޟt܋�6�nz�q3���eׄl�$��8>�#�q�XJ���g��!/�Ԛ��y���3�f6�&�Z�M3�Vz����
1�
/��eR��п�Tv5����>�Ēږ��� C#_�hg8�?����u�ʋ�j� v�I&��5�z�پ��줒_�[��xPw<W �a��|��ȩ?j4�9����QǙ@�ө��[���ִo��n�w?k*J�t(��C_�b3=���g�9�:�Y��ՓV��@�NBG��������G��3z5 K���j�i���q�`=�`RO!_����$At%��s�J}$�M&�Y1K�Ut�Q��<<��N=�"�� �ha���������\���4����"�������:R1�#���]�m�^j;]m8�����JI^�i�[��Ƶ1#&Tf~���q�8XY��s�8���Y��m �V�����I�#X�k}�7�V�{�/�����R�pD{�T/����QQam���%K��㲞	��N�b�/t��ݾ;t�Yu�@�%��K\ccS����蝍���4G��Z��#q]c��ᱮ?�����u��]��?�:��Uq�o���p�?6qL4&a="M���?whcY�.�#��L�^�V��Ь�uzo��#�.P�Q���ؾ�ɻ
��Aܫ�Tyz��!_�~�Gbc�X�j�-پDfY�����p.��!W�Pb�r4Vw��Aij"CU��A�Fvм����<�x�Ou���Y+���G���`f.ɠ��}7��0&��[O5��G\/M���m�� ��;�1L�\���Z8�P���fu�!�f�+������_��&��P�!{�yY}�<�ǻ)�l� ��>E{3G�����;�����tOZ$@�I�wkY�!����Ĺj����[��y8������\E���|W��͂ Nf��\��<��a���/��𪸔�k1�C�h�03J�X/E��ʾ��V��3�����\� y�R+�>��H�U��Ē����uh��c��)��^�d
���ϓ(޷��F��ּ� �4v{�V�^Y߳�]�~~C�D*�8.H.W		�:J�	��䳛П]L"�#��ګ��|C2��0I b2���@���r�II�f4�Bz�[�3��5����OVN1����u-�׭�bL�Q��L��tB�4PA�b/�!Y*�:��j�<�(�څ��
����N�.H�k���{@1����y*l����G�t��F����39�����\����-���K�*�G�ǁ ;��.��Ծ|nF�lWv��z�|�=���L�㋞�PE!� �[w�\-I�� ��Ju�:l)�e����f�Oad��86�|@�����@�a�`T��O䴢׶�b��Eb>�*"v��Ӄ@NT��9X�ZL��j�=lYx�PV�9�i�i �IPg�pO��P�S�ڹ�����R�iA��AQ#�ɩ^[B��*L��6�����$�Y��o*�-]�I�w'�N.��,oM=f�섍b��F��F��F�f��6��O 3m�\I:��1k��L�����P��ɱ�tU����;�"c8"�3����Hl����зd��.�T}"�Z
s�8�
�0��|}K���J�i�j���h��mG����,"�ٓ���:��s_�0B��*��ZF���K�kpC}��^/��r�� �Fv�/���"�_�ϚUf~��������;bFp���BF�½�L�=�}���T�_�4��6����1>Q|�~C����=���s�11���܁�]y�މAZ���g
�N�H?�Az�"����Hݼzgv�����6]�X�^U�B����b�ڮ[�ҽs�x���WUY�v����:��X�+�$i�Y)�����C �y���G��@�/�.{D�=uc�5�2�(���'g���6(��b��߽gPy.W.G�~~��vj�K��[�P��/��%90�@g�=|C��<��fp��j6Ah*=W�t�Oȳ��u@�c*_=tr�{(É�~8o.u�!�h��+٣^[^�mѾ�<�^��EЗh�pq��n�~i����1o6m\8&��[�cִ~`�-3�"U�	�����lm�=Z�D���A&��rۜl����99��b&?K�w���xmM4�R@��mdc���or���L̊��5�Zx����Қ���9z��5�;Ҍ��`�j�oA��N��y妦�D���p[YL��p�
���Q�\���t��5��1���8!hV�Jt�r������wU�u�:pi��?�HJs�Ȃ�ԓ|~��p)s�@,��`-N=�yf}���
���A��7H����]���0��p彘�9U�HT�h3^��H���̽�f|���N���r��
rS��?GKb��j�9�_��XUW�20���E� !N�9���4~����\�Um5Z`���b�Z�I«��3�J� М��/�®�����U/�*��,�]���Z����Eݴ=:�#��5��Z'�s,�w�����I�Rj�$Vîz�.a����;-d�V���t
��bD���(�a$I�lջ��?aD2Q9�J����n���*WuW3����H*�����Z-S體�HL)��6�'�\����Sw\�X��ԙ�iӟ���m�N����x�_�����[��<�S�.�qVe��h�\���sH�PS��>"��W`��Zv~�ȱ<>�#�R��b�'�2q&�䴣�`a��+�\@�7H_nT� �V�(��%e!��K}��V�E��O�C>�����ˮy�5[���-#У�B �T�L�qQ���0�z�@Zs;o�ǈ������	_�闧^A��\�k�������6n�-��8��ü�Y�"������`BG�/f} ��ҿ篼�2�3���6���D��?C�{�ђ���Ԝix���Q�U��'"�#����]�e9� 幌M�-snW<^�?���o|o���o)��n��-�,M�9���ZԵ�k��z��v�P���M�H�,�Ejs<�J��L�q"��E�{�ϮO��IG7�sm�rc+O������5���m&���Z�(���o���@8E��f�R\=�?�vѽ�\=:l�bЊ���T��)Ԉ�N��9=Ađ�~a�<wf�!qi����n�Py�r�N���M߈Iix[�|�D�|uI���p8��\�F���@#����r�O���P��g�F9U��4���n�S�¤~0����w�0o:Oژґ���ڒ��������֦��-*�y�@Hݳ�(oC^�F9k,�O�f�z6��ǓH]���oŏX�\����_E;6$�F�-��U,���_hd73)}�RK��8�l���Y^ƥL��3�$�ν�A�����A�@d���r������ཕG�t��ט�sf���Iz�o�g��[iV���^m4����k�ܾ�v��|O��S�SB\8�w�[ E�̪LH�7Q�����w���cp��|R�E�ԳD7�\V�M��Q�ֲ�'%.Q}�Q��?Vw���Ա��%lh����z���I�ħ�:Ir��Q9�,E���oY��J��')v�Z�����vm�����M�(;)�'X���#0ԥ Ul� �5���,L����e,���up+9xhS��#�u��&�-(�]�M'8$Jl�8 �lM������4��l�c����70��=�sq�����uO&x�W[�W����ۧL�hG�`� @j}�=*��^$e^�FT~Uc�7�����c�5e�|HU4#��惨�4��j���2sd��K��_H�5��`�����J�&R�m����sU42��̎tۗh�͹7-�;��8�C���������8�� 8#.��֕�O�CZ�qMI�v����ZÇpDS�!�C4��P
t��=]���{�2Kj7���O��J"C��b=�#���5�t/��B�jA����M��U�TX��X2�
ԑ��I 
��`�ym��Wv�Yf`ޜI�w�_p�>��f�BL�ڏ�0�Y�Q}{e�n���}��)mB�5X�����z����!'��>����wr�U�=&�M.V��R�Dk��酯�ہ	詒� gșZ [_m������zJO��7��@`n�"�@P���嫲!�ޫp;�����P��)��t}\}�����#��o6��bB'����dT_���OQ3Z�V3��mtô����c1X�������gf!�����v��z�<,�����u.b�}���P!S�6�ՙ�X��Wl�1��7Iϕ�0��vk�ڄO�g��w�a/��6u*> N�!���)������=�4��f��qJ��(�֛&����p�'���װ��7����H=\nDX��^��&,�[�h%:8�}h+�lZ�r�
��N�k���D޺��T�pgQ"�_��3�>�v�� j�b[p�^�3�M��բ���˫�m�>U�eN�����QX�+gV�Ey��7�n"�Y�^0�L�*�-b-c���ʡ�!��q��ݶ��.|��	�',�H�Ig���,tEn�&6�#8�s��,���5��Ȣ�.�������i� A��-Q��)�Z�����aE7Gޟ��?��uY�G@W���)���V��V�~�r[u�h[|dT����Q��͡�2��rc��w�8H�e��U����:I��Gք��1����˨d���6n����X���űM�sU �+����h//"+��l=K��Wzbm��=~_퇞�/��R L���2*��*+��e�'��{�'��Ӓ��nI0����q���S�XPɱ�J�����\�b�=�"�"��]�q�$(�����d3��>`�G�=�ld%7�_�kzu�b�j�4���9
r4�����o���,���K��J��#%-�~/jl���	�f;�R[�=�`��81'���YsMݸA�&QҢ�;̆%/AR`�yۧ���l�ȵ��ut�-�/a�G����T��w�$�=Z�Y�'��fPW��\�J�*�)�+>��_e��a�Iɧ/��	�D�'JQ�R��( <���n���d���u|s��f����S��,�cN�x�Vޥuܽ���M}���-�x p�d�)"5���|�i�)��k=��32]�=R�oѝ��je�|Z�S������m�HR�бbvAK�]����Q�"o�Ӳ=��)�<�O�x�T&�����=�ё7��2�ͭ�.h%�@
����b�.�4ļ���Z�vD��1���vƦ�l�t�q�C�{g�`2i�Cg���$���3޶���p�1agZ���?(pf<r&Oa�8*�|���	�"?n^L���Z��Q� a�����d����.�Ϸ>�\/hbр�5Z���4|��v�i�y?X�c?�Y�q��+G�+�O���nNX�P<����Á�Q.�է���)���Qӌ(��[2�z{f��$�,�����e����ճ���矙�҅h#���
���`�o8��� ϩVk��F���|6E��4�k��_����\�<j��y��&Rg<�����PCč1����;��aβN��A���C�w{8 ���w�8�
���=f�{-��0�~�M�W@��n��\�`��qo*ڣ��v@��S�2���4�[������4���Y�v�b.���$�{������VȆ�Ǫ@P,��8]�}ѕ1��Ǹ] -��G�����č,��o�[I�C�.��$Ϳ������tK�ى\�&��b��u9}�$/HՅ�B	�W7�7}U7}>G���X�[c�����<Ljt��0�&2����5q,�5�P�F��6V7q�c�d�Ȼ���v�aM��_��W�oVk#ƈ��P�%��4��,Z2&�2߀���ؒ0���CdM
N���Iw��b�����E�a>Ŗg�*V$����Z�M��t-ۨ{��3��j�u��[$�� Cp�~�!"x,�I0]��i)o֔}����!��SIJ��'�KQBqk�R��݇��ȇ��Or��e��$^�τM|���j��G�\tI�DoR�v\aPho Bɉ�(�&�"�8`w�gR9�;���#ِ�ZT�H'��P͹m�{�5i�1�a���mDl�<'!����u���M gPq�F���b׺῞h����,����B5!$6��/X�Q#;�Y����:%ΈJ�b7�o�W��*d����f�$R���CU�_^"B�# �F�D	}=p��-�!����:�@�D��q�DOɀ����J���q��(3��U??v��ɴ�G��l|��	�߼��xI�J�c�U�p|]�7Jy���Qypv4ٱ�u�l�h�ǎK�_� ����2��e� c�a:�D8���!Mfm�F7`��0
��e��7O�h��y�Ŋj�r�W���#�AP-����N��?��t'LՌ%y�0R�M���!i0�[�6�m�Җ{P	��U��oH�Ms�t뢏m�����b˩ӽO|�?1��%O��
s�9gBO��g#˜��G�	��.0�7R�����.. �<��TM�s#R�my���)[�~
�&��lw<J	8�����&8"��}��W+5s�m�]�Ħ�<��L���:HSf�J,�y4�@oI���@����?RfC�ͣ��J�)	��	ģ֨��0� �Pi���o����m�3\|
��~<�{b�$�h^����`���7��%Wx��qA]��E�v0�J`��4~�״�N������E��c�M+G|�N�ωUDf��Ʋ����תF���z�ʸ΀Ka�kB�S9��k��	��GE�@G���"��k����n�U}C�����?�x�]Y�d>���8�f�c~q������oj�Ɔ�"\�EH~�h�G�:��LR~6�w�?H��o�u�Ѯ[�43���X�L������:d��H׌ɛ��}{�;C�g4����my��4Z�>�#U%���� A�(u�"	C>�Z�A���,֙<
B���W���P��^j���zutK�K�7����eJ}�x�2�b���ֺ�d!�Ϫf���v��܃,�9q���5o$�W�������A���%?Q]B[m����͝Y|(�ǌ�6�� �� �?rq=��S�yI�EO��1�
���$Gq��F%*��;1Lr#� C�Ƿv�0���܇�fmx �o��pl��
�e��4����g�su-gpգ�F�ݏ�J��� ���)x��r�U�J(,ߋih�j��%�6.̈́�q��&�-�*H���#��;S�-��7|/�^�( �V�n9��:^)���gF�:0��!����	�/|�@�t�e�h���D$Ӣ��I�X���0�_	:0z�c�����/����C3�
��+�O#��i@g6��i�L�^hw��v4���	*@LS;'�H��Vİ�w�ʖwPȽ!$M`�򖗲L�@�bs��)�d����'"6w?q��p�j��X���v�S$�.�{F��lȳ:����C.su�[V=��{gu��v�n��K}F�xys�r�"�v{��s���P��m*�F3���j(�MjChl��*�N=]��N��p�+�U9�U��bm�٧$5�x��}Z�Ky�RNn�+F;�����\댘mڂ0Q�_7���r�m<ᵰ<��L�A���	�*��7Fԧ�pӄ�?�*~}��D���������:�B$͸��@9p��d1�>	j���XD�4`O�
%Yc�<��)vg��q�@m���T�����i�m���wx��=�i]��X��0�����xx��� +.4�B_�gM����eJ4*t���WS�AR�<�b�6�7����ٰ7�/Y` l��1�Ka��-�J�΃�OXM|$��u��샿a��^'8����d��������8��Q4*�Ԛ��R�.ʛ�/�05l׭	;D�v�r�8����f�ꆤP���_\�Ry$���ܖ�D:�Q�D=��=O��R�A���@�kaO��r+�����z���,�8t���>-)a�{���K���$	X�7��ꍊ{+�&q<q�a�!?^�k���wa��ae����詂�
4i5��u�D	�Ld�ŷ�w�t�1�E>�r{>�7D1j�ѐ1��M�ˋ��Η��5�o#2щ:5��}3�EW�8�o.MV�;򁾃���5�Sn,�F��dp�q&UU��˧
V%Q��15�&v����z☄�9eE�:�?�I�b	�E��y�hwȅ/a�{�cn���G�Z�A/�*��#���ѿkoo��ko���X���*Z�ed�1|~������QD������Go��cM"�Y� DO^�e{~��e\��iE�g��AWN����K��P�ܗa�_8R��g���Q�*~P�x�Ŀ�;e���n"#�SWV~n��J%���6]�fh[P ��Z�Çʻb���+���D�.�3��OC�1�R��rv����;��ɿ�����RNN8l3�t���PH�����L���cJ\��@����9'/\�����o�`�}2���Z��0�x}_�Cm֤�iWg��۽���\��p79[M�7�#����RYx��5vоy�w3ε��Ȫd:ͅ���Zx���f"��u�j@-�*�G.PW"���olv��
 �E�I���.g砋��(`���J�#�\	�)�����H�,�5�CB)��9�Q���]Hc��C�����G�W��i��ZBk��Rw�O1��Y2�F���(�7�ҝ��lb����%����r;�MRl��N/ڨS�a�t��Z>��Q���Aߦ-h��gsH������Lw��������:A�� <A��N#y�ׇ�r��ĲRnKI�]������y�t=���2D���Bj��v��^���z:m��j�I��VPA�@ms����O|���~���7^���݂Ѵ���0dP����f_G,ǅyg��%�=�+ 7��F���L�rJ��<9dV��)�3��FqS�O��4W������7E�hQ^�Kjź�u�Y���P4�0�}ag+׿�	zy�t2�?�Bu\0|܋�5Fb����A��	R�c�*�^U��$mP� �|kru���U�:��eKv�2�c_t\Y�1��i�=�$��N#|� 	�E���>��P���m]���i+�"�]�T��˲rH%J�1ǅ��["X�H�.�ަ�L��{��Θ�!�_k�d&K���@��S�MВԙ/����������_�Zl1�n
+���*��}dVw�RF"ESG�}�?v�zA�vg�ͤ���|%�, ����ޡ��ᗶ(��ݓ��Z��;�U�r?m}�,,�5�Q�V���ǐ`�K��/���<ś������Rm�xp��Y]���wYc��YG2N�'M��h�~%}*͈~�m�V��v�r�yG/��J��2$&E��F����_���ݧ�J�3�t�܊�O#�����H�%�A!&|,��:`�"��)���:D^L��%�����hn�YݣY��ux�wSk�����
��{�U�7����do�"r.����G���������P�8Md��F[T�;��U�iˉ����$&����}�,��DDp�$J�G�������B�\xrUzln/�D��~�m�R�����T�M2�@x�ط���:��1Y���r��c��@Ў��6_u�L{�^���y$!/Qu��ݼ5��M�o=����։h͙^+[W�,/pq;
l0�}oۈ�ۊ���g�2�ŏ�b��2h�\c!�FdJ�Z?��m�\���K���j�'�3�4\ѫ�F��x�?���p�+'�x��w��:?��u��zʪO����`��d_���o��?�ﱩ~K���~F����z�+1kp2�Gg��qW'�vy�;�\=�1����%~��d��������Ng����+�%`�:7FG	ɠa�	C9����]��t�4#�26�<�v�����*������!͕�vܑ3���Vz�F<-�V��<�(�������m|�h#����q� ����STwdu���A�dD����~���i�P��a�.q�x_o���r98�*�	^MlyK����%�; 1�l�<G%�� �^Cmf��u�����p5#{a��)���l|��C�8�,<p	��g�*�!+V�р� ܵN�}��`�2lP��D�C�`���h��PV����1@��G�G�P����o4�؜��f�Byd�<�R#.B�<H�A�����G阮�����]a�4�U�e�T����͡K7����]s+V͉��%T� �]���k��nU��~-)�q~ph�����^, Q�:�����c�ı��4l�"Z��F��`)E�{{LC_����-���^,f��:I�`���J�W�G�J���O�y�"[S��)��+A?DWR�IK����)��^?s/�:%���92� ; ��$X. }�Ah|�hd~7��G�?�?s�h1��<���a� P�o_qdY}Ik��
�ђ���S\�,����(Q�n���h�P������,���B���޶�N4��4nJ���f�K��v݇g���v�������iLO���\���-��@oE�˦~j#ơ�8�S��^��řR	�:�;VdЃ��A|�T��������lWP��Q�+�����s�^/������a)|^J+	'z�k@�]��Tyk�@�ƒ�����OY�^3�p�P��7u�\a�UwT���m�̈Ϧ�������BQF�q��0]��dR��*�z2;������l�z��Һ��1~�}d&M3Hf�+B"�ѾÓ�oR�a2�s"e�K6�>��A	�7 UB}Z����м!%�^��R��!~$	7�ɗ�[���R��V�#��ع-#b}���6����_V������i�..�9@��DKGI����s4΍rl���]�￱0�svk}WQ�(����5����8�k�&"���Hq�!�{��+�2Ԣ��[4�(u�?qD���Hx5~�ԷA*Z�n"x�!0�[��bl}�Ď���gj��B��I�n;|��ͥsTEm&�U���=�ǆb�z?Y���&^�p�����Я��bܸ�0>~X��Т&�4D�N%lUtxP��� q�D��JAm�^���9g}V5p��<�P&���cm�X�J�?�g�͑�X�=T�_ժ'��e��d�j����A��nI���,�E�Z>}	��D��W�Z��F�B�|��n�sQ�r���;|�әn˘1���X��/~E��T���up�0��Ɩ�|�36�(���ܙ�>=�^ ��2�4V����$@��`�B���@6W�'�8h�^mb	X��A�L`�Oh
ڷxT����#�������Mr �Q�pV��l&p�b��%�&���jxl�mTC�~����'5�V)�F_d���Nö�����1'�gs"�m�x�@�-�*�������Kj��$��ߓ	�(����E��&�{t�_HPW$�nE�uA3�c2��Iz+��_�G�t4��>ˇ��y��;�,꟤j����P����H	&�(�V�z
���=nvߚhKj��<VB�|��azg�g<r$V.���m$;�3�!�/1 ��F�5Q:�4���1 ���JTa�	�?|�!�s�E��fN`B�9G~ߣc}�;6�1`��M�˰!c:��)�T��R���Utg�7�B�C���^[�cMA�Gd٩��	8m#"��q�	� wS���<*��>%�7�&5sNLh�?y�W� `�h%�#j�Qf����R��s��v�dX��K�v�o���F�]�՞!�OOl@����Ƌ!ZAXD�#'��0KX����U]jH��Ad��&vvB����SXB�WUN�0c�zw����+��*��g
�F)�顇�l�^gh/8����>��*�C����3�՘��O�l�h��)ƞ�Ľa��U@<�l?gD��@u�����b�U�#��W��a��x�>%���*֋f9(c�2���pyA�l������gB�C��1�?O1TjH}�������WPi��9�~��Ҳ�ɠ�\�Y�?�-����~iO��.��S�`������S���w�^!G�Q�^�������;;��j��>K��.2�x6]��=�E{#͞g��DB�͝tIEK͞ۣ0�� �宜@��T��$�ٕ�&���ŔY`�� �:/x�� !��-�X�{?�%X�y��},U��N��&�����i�[�ݲ�����a�+-��q�«�T�
�8�����~g�&��s|�
ϑ�S�[t[��u5� ,i h������5����!�q�@�VuyxYY��q]��
x����S<oh��c=�1�];�p�零jb'X���"v�/+_�<�ﬥ��c�i�U��YSC�38V�\&Ay��@˚E�Q�SPvX����'�d���]�B�[���ˣ�2Y�}D���,���88�S���P���̢�s8�]	:F��y�7��|�Ń0���p";@FP�㋶��p��ϐ,��xB+����[#fW����vu�!�j)���D�ڇ|w����>���e��MH2N]7t�����JU�B����)����#��Y&��]���}=���p6���݇�*�%�|2�A�sU��^;=d�ޕJ��7I��b���S�����[��(O<��]�0*��Hl�^������:��2�?�b9���
��&�>Mz^Z�v#t-H ��A�0�ч�O���#4��4�xM^"�?7q������Ji>�^Rz�Ĵ��
���zZ��+�i~��[�ʳ���ՂԵ��q���+p��g-�_���%kDhL,A����ď��q�O���S�����]��6s��A4�U�N��Ͱ�؊���E q�� 8���_�W	Q��6�&Y�G��|q_�$�L`K���8�F"����v��D�hG&�1�E�Z�	�娘?{60��m�;{�Ɲ1���NJ�o8���e���R�eż}[�?-��";�1ni���t}�Ԗ����{��!��sh�
�cMd���|���ި֪���lq�"X�- �H���J~�v-�F��|I}nj�@Iv���l¬ge#"Q����m�+u"��	�yrI4�\��.��_�1g~�I��#���F\�qm`�"m�8�8��ċ>���jLCm݆4�����j�i��s/�4�E�u�9��H-���V�c-�~H! ��;���~�َj"b��^�P&�)r�&�xD���f���#�ETu�o�"-I�b��u�ysz����*��x�?/�V]�f]o�H�V^�@g6�K�I�G�/�4_	�K�V�l�4�h��t�/~�6��C!����?�+&�~.��ү�=�	�pji�)o)=����r��?v��cGO�ք ͱ��8�o挐��*�z�z�=�x������,��y�0��徑������0ry�|�����ڼ�`
V�7����o˔:NUl���_��=����NpX��;ʟ4_L������X
!��3���n0��mZ�ҔVa�>��JtQ��(�A�͇����a�.���C���4F�WJG^�,�������h�dhw㊹{e��������D~%`?���=]�Һ�����}/��,�"��?�M�Vh�wg�ڴ7�Mv�QS�[�0�t �	����HB�4��4lY��Zhj٠��-%/ib2�0g��r�A��D���ͮ�޷мpmS����7�?��q5}��69o��,��|n+q�y�A�7��Ҹ��>3�����H�Oj�3M�����V@��:��;L��PR��ɧ�V�L�F[1ߕ��!���f�9��
Fv�u����O�?�L��
��k�U��iAr��1O'�����`�;��sؾ m��g�(�*��n���D��w�'���n:2��?@�c���Gg8�2)C9��F+������=�x�1��R���w�J�����F�Pch�̆�b��>zηPkr�d�С�2G)�2���ݩ͆z�l �F�M��)n�nR_�a����]�A{�']�:�P�H�)6����W��a���ɩP�O�������c�����(�+U�����'?=y�ȸ��dC����Y��S�w��/��̤Z�l>R�ڦ� �#h��Y&�)��W�h�摋�D���'��!�d[���ҀF6\C����|��~-�Ņ��π10
p<���;}˦'͟�<���e��g1=NC�c�Ҿ!�xi�H�v<��B.JKVA
��H�\+��6B4V�Pƪ� ?}��}aX�$��v��k`C�I��tk��!�9�T�bRa���Y,fp�L����)î�����|��F5:�?������������Ny+Ɉ���1,�m놮n���N B��X9;�ɭZ�t����p��i��ڭ���8{_�\ͤs��c1VO.J��6����(�Bi�2W�N>���^wF��J�
�c�X�Ѳ�����+�߻�T7zA�
h���-M�E1���y��y�B֒CN�)dœ�M(B)��c�*�/��$��IǺ���@�*so34.4�3V��9��t���ڦ�{�0�)���Jڟ�6���_ǊD=�O��j�|��RuJz\p�����u	��=T%%cx���X���8�dř�ײ4��([]�-Y��7/��51���va6z ���1����(Xh�ղ^,��oN�erǇ��p4�~R]`Ƅ�������b���p6��L�fU�e]e��F ��]&�h]}�'"�`I(��ʶ&��n�r��"+�ߊ�<��G6�V\��Ur�� �-`h�����YZ�W��)�&��dq�mt(c�nUx�$�Z�P�M���t�Nz��>� ��O�^qv�q�	�2a�0T*dŽ��0�fnt�uX�*�V٭�K:�� g�~�8À�����p��Dja,�㎣'VwTPڧ�x<�Xl��/�"�q�����m�0�	��r��*��.I�1WOe�����OU4a�xnY�W�|��y4+Ekx{��#�y~�4v����g�Ztl��`���h�Kr\�(�c�[�_�ى$���[ƭ�JB�C�\��w(*�i��5(`�
�6����G�ŀ���B5��c�eǙ�N�߽p�|n"n��k!����\���e����4O)k�(�#�~p�~�¾9=qGŇ���8�h�g��G�g`3$u��5���m�M�UD�0�ꠍ J���Á�>�ޓ-v_��۶"f�]�%��~15+9,�BtPq���.�;E����T2�O�u�b�
��н�
�g%��+-�7M�Q|t�$]�?q����г�1�ʣ����` ����4���t�Q��L���q��ތ�fTgסʏnߖ򌧛�wY��u%oZZ�-�������@f��;'�B� _\>�n�AR�p]
c�#��ի3\el��������9jo~�&�ׅÌ��;�rô�����vq�UJ����It��5�{��ۚ��ǃQ���:Ee�]M`�G|����`ԡ/��Cć.���Y�>"�����k+E=0VJ]rH��I[�� W!O�c�b��
6�WB*t�r{P D4D�*��p<v
3�˫pi�Q�%e7�n�>��
7��h�lS�"����189%dL�,�d����Z�Znۮ�`V�P*�����>�+LS,�4�̴�b��D���64g�h)(�8o��F--��\����8AU�a��-¡�_����%�)�ެ���	���W�^����(ʆ]�g�v]���x�8ճ4��[�Z�@���a�R�>�,i��$ uS������ ?�&H<����҂?�+���������x��_���r+Q�#���*3�z"��]��-��Lr�������槤�����`��=�4U���;��|���ۿ�g3��#�Iӡ�
�Y���5��{������������/%D8mm�,�Z�e�Vhx56Sw�R�,3; u�_�w�ZF,lGh��n�$|�n�ɒ�0�:Z{�M��g�|������p�e���&hk�̤�V�1�\�t�#i3��v$ƨhLg�:��<l��@��r�נ��Y�y˼,>��5�~��M���R�ǥ��*jQ[͙�~'�|�v[��c؞^&E�daw�����b�@�Y����0N�z��B�`Fa|tQ���#K{5C�
��l��`��6Q��"��`	�d��l)"��(F׿�]����!��9>�7�H��7e�/ҡ�h��	���	[긠/� 	�~T����p�'�qf�B ��"���R ���.�ܞ�7�@�HB��s���殌��a=nu��������%��B��EX�V�2`w�#�]-
��X�C��v����BB���la}�F�N@RU��R����23A�=F� �+�;rS��b' 
?����g��	��3n/X{���v �B�1ȭ���eO�$N�$�� ��X�����yq�L&=�X5�������UZ�܃0X��g��'��.�c�o�f?L�w�9̛i_J���B��=>�_�H3��"�_Jd�L<�U�Ыx{;�

&@�f>�O󻾼(.�c@,|��:D :�뢥v�Qb�����&��i�(����pw����f�64�K�֜�y��V�Bg=��{��������C�����u�Z'Ɏ�y�$!�yP�P_;-��33�1U�'V�l�>s��ΐ�ݖ�����Ѡ��^������	���cX���P� Z0��Å� !�˒���vLܝM�M����^��5�/o��^��kQޭ���4cv�9).�7œ����hPwQ��v����I�I0�+*ڬW�N�#����=Ùgw~]_��$���Pӊo<����b#?6(�rtɤ�(��ĉ�J���f�ow�"�'�� ��YţgZ�K*�H�E��M僓
��|=��}X-��c�����:�7x
 �W�i� &G���ZG<�Xi����=A�"d%�^B��,�n3�eZt�t�;Gg��a��-e"�I��<(-<�\e�f<QPdjUŁ�{�n壤����a�N3�m !<~uV)�5|�	Y9t5�DO��֠�i�;�O�PM����W��Z]�ƾ��,	ķ�x��3��V1b�� ^��.�o�h��ؔY��/B�F0��O�1;�qC�@G(**ɬx������<�0n�fZ����ýH\��q���S��c�������P���:(LՐ��1����FB�?����n
v�=����t�h��j�6|�zf�yw��6��qaNNZ6�8 C�Z�y6��ѡ��b�Ĵ�H�Ḹ�c��R��sm��^�og|�P�%��J5`
$�ڬ5�=��̎P =����d����ck�K�/cЁ����rQv�֪^���x*�O���5\�5���}�P�zc?EM�0��|3Q�{)o��'��/L�U���
�B���d��ʶ��4V�ኃn�nW�����nI���{�JѴ	���U�{�p@6�b�Qݨ���?�'�f
�;1�}�UuG�B<!9 ��1��N�m�%��Ԕ0�Vi{�#�\Q�Ftǉ|��6�j|FD)�����M��n�֥M��ӭJ	-h��cI,��Mx�yQ�`&��y�v.Ls�i� ^1O�e���� �!hmy ��b�Zԅ�U
��:��'%u������'�	�!�;�1�ƢZIr�,�!�Tt�-96&��#��G�bnjF�6��ڗ电AN^��\�{ض�n�sNV'�S�yV�=��J��B�OBb��`����z5��1�J�bҤvfus���,�b�U(�臛X�y p~��.�$4�fK� #�m�Q���Xد���"�3wt�u=��
8�LRdٙ���v"L~�����D�Ϳ��_�0	εz�v��'1v�W��!�F��*-p�D������`.�F`j� 7烌D4ހ�Me��ԏ!t��{,�O#0��l�&��p}��_���'y�ui�'h(���g9�Uaܰ����T�;�po�n���K)��|
�6)��DV��A�0_���O �,�M�f,&�>���/�s$�%�Y.~��Ԃ�F3(�ɋ�v����4�0q�H���0���"�Y5��E�O�t�<�21�~y��~��%4�%��Dl�����M��������U�/��]���8�l�>�"<	��T�(�(�j�p"hJxi��n��%���¬�R��^z�m����P�G��IcM��$�$z���GҶiSo �$&G7ղi��`�(|>����]$�{�Gum_���mU�YG�F땔n�F�K�4����7�Y���Hy�������\�d~sU�ϰlbʻ�M3�:96�J%}�|P���K� t�m�k���Օ\OBĘ�Q��0�Aj�ջ?�I�ߢ�+_Ϫ w(�l�aiT.|�H�����j:6]qzu��kS�]i�SrN����r����r�#��v�I	@{w���t�_U0l��3���j/b�MX5G=�	\�^��0O�Fd���8��s{6���ro��%�7�qS�n������}�҃0+C������/,�YA,dbƎ���p���� �]h	M��\�����Re�����,C���K۰���JY� ���m��Jɰ��ȧ\5I�F�'5��]�����]:�3�^�`��~�!�B#��Gƣ��V�YM�xXes�T��m��-���Ё0��D�H ��*#.$Ծ�^����;�R�2\3�͋d~O�z�H����B���s[5H@��	�na�r߆8�� ��o?StT�`��:�x^�y�����_4hH�-"W����ɀ'^<�}B(5�|si?��� �s!YN0uh�v�O%�,iz���s�t�ַ�+&H.�	h�%��I4� ۾��El���@ QaCoH��jlf��6k1]�pH�A�Ҳ�rZp%��֞�@�6R�9h�nӚ�����^�v
��2\��C~L��Gg9�A0���jC��������9���Vb��Lg���j&�l���'�����?��#s�.���M�izI��<xG�9d�5��u!ƈ��A8�uu ����.�I�CS3��%2�rON2���R�Cx�l���l)%1ZxW�,
�<�����B��qW���$V�»�+WH�$�X@9����z5D����!�3,��Rl@����x}Jt�c��Ems�v,J^� ���E� |�A\�(�|��Ch��4�:��ܤV�Ե�\�oN��A� xU$H�t�������S_k�����6�.1�D��]����yO�|����EnM�(w�g$Z�	t(=���|jy �b}Q�F8D4��k��H筱��v�Yyp��~o��*4�=����=O�����ϔ�����/�_�c�v;� 	�CT��L�|�e9����cL������7:�5�1���~�۳Ե�����F��4Yۗ�)����	 ���^��d�͉���IC[Cz����.�b��_3N��ug��[��@�V��ppL�TC)��Y���}�R�.��d|�+��,�X
�w�C=_�\���q~I9B^o!1\:�(����Z�F���5*��v;�S�N�Hd��C"�-�ԫ��<+�U���Z'�����ʝ�=�ǫkiJ�<�Z�zoP(@��߫��㈬T���$��7&رi8�3�;�Q+��y������F`tS�=��~)͐\ f����UN.*f���o����U�Q�ˇ_Ϊ���2�c�)Ndu���@�$���:���5g�w-���0�I�΋q����Ϸ���Ma�%j���6�.�䥏D�<a�x�L�f��lC;<"���C>q���������Z#H�ل��G*��8������@�|�w�>(ŵ�ބ�ZU�Hw9}�[9�g�r>DuDl�7^�664�Ϊnb�Jǈ�3B�SL�U�2���X�U � Q�	i��I��ZZJ�1��6> n+�nAr"��(,D�	�`c�/<@�xg��%��qZ�5�ץ��`}��\#����{�F���,�ł�ӱ�{CG��"=�X��!E"x��~_.��oz��q�-��aA��S�ϭ*���������o��/ )��¼p���S3�W��vD$.���|NQU�=	?�Q�X�BJǺwu����!�����D7uCb]�yHt���B1������rn.Ñ�z�x0<��`�7�;�ԵAP��o��_ҼJe&p�ӞMв����gv���3���_��x������}@���˥��~9����E�Fݟq�Xkg�@[�}� a���%��c7�l/C�|[�n��L��wh5z�}��'-"�9}?�)����΁��|J���Q�?Пr�p���V�Vc��U�aXsU����@���ʘ�0ў9�Q�ֆ��GNU��	Qe�}���l-�vu�����@ �ܯ��X�Y����m���Ύ櫯�}���ƶ�0QCRf�s����ːF�*4FS�<Z�X��N���\�iW�U�y�+,y�*{��Z�C��a0��P�s"�㑑�?�}��@�Gx�����T:�H�=�������R%Oj'����@>�BP�ݏ�-	�j��ݩ>\���v���#G�{O��s�~�I\J]��?��D��T���&`��8�6�Д�`�����O���C��7 ��I���-�ь!�q�6,if?���V��U��Sx�#��-#?9�Gئ��%-�K6N��	��M�6��r>��0�X�\	6� x,R18{����ca��������$�~H�C����o�ke������C��U/-�Bg-��=��#p���e.=�L�3!K��{]1��xA�Źjیh�L�d�ȉB�U�t=�3?p�/�/r�.Z\~W�b���9YBS&gT�w���H[��>�O�Y�1��M`Q��اH��cj�`���kjL�k`���:
���1����������i h5P�3o��i���H����G�b��k1��������ʵ1�!
�%r7�V�7T�$�N��nц5�_O��������[�x�{'�1�a{�5�>�5�5=R�7��Φ���Ce��&gu��@8չ� �O�}�#���ޡIzj���9:�)u��r�ڭ�����!|j��1��φ���e���� +n#���� ({'c�@��Zǖr�gBG�o%����
�����p p�S/��q�
]���r��2+��!`y�~����\t�)PO�����j�m�M����#<,
��v+l� 뜉��w�*�%�M�����2�-��@`ܒ�<�^��_;��qv'ei��(��*�X��NT2o��k�{�.�^}��V ��(x���J���}u�vhՌ��"��/����VK����nK6piIl��i��86	�����<l.ӗf�sj������LV3w0&�A��9dk��.uU"��R��R��F���I7@�%E�ﰞ�9���=(�?�+�T�_T&n�0�$���T��"�Xk6�?�72���('7����D�4^���ԉ���a��m"��o���?֛�&��&��-�{)Z�P�䔠T�@"�=��� *���S�߾��`?u��-��n���h� 0R��	��@)�:���r��L���?u��"�!!�����S��ﾴd��)BU�� 	oK�������>�q�󍓉�8��&��TPTz�t1r�#M��-��q����R�s��6�YaT���D�>�W���Ӫ}=P���/��z�H)런�;�\[Sp��bp�Y�c��ے8��x�|�@�%��H�?�"oN%Y�/���oq��c-��*�N�)����	z��IJqYQ�����c��(y���!&��6�K�vdv�EJ��cZw��3>�z�߃�?@��n��x�]4M��i��O����j÷�g� ��i��"C�3n�{v괵��^!h-j�h�4aj�XP�0���:�#ឝ붟w7�͋�u�Y&UPVn��v��iN�S��
V�P>n�*��(d�?�	>ΑA��1_^���ϫ������I�����*:a��|$��M�y�D��R��v>UJc�0MNj����O9��P"V8rƘ�p�L0�fm�_�j�f��UI���kΔ���^;�WTq%���S�*��ү+<v���i�M���d�˞pY`��X�>�}]�`�K@�H$+������
N������S�ޱ��؉&@���)BY��X�J�����8+��P��f+�C�A�HA�+ƅ����4�е��숍}��tm����b�'��6�&��&���o���ٍ�}$D�YP��xO�����4����K7�$G��}��*|�8S��4ΝZ�M?�>��Mu*/�:�4������O�e�7�B�/�q`��B��ϖ�����z Y���I� z��xv�~Ĺ�-o�34[��$���������2�S���)�Y���jӶ�b����^�t��^�ӡ�ȹ�yB���o�s��Q��[Jy�RR��xe�)cf4�w=�	���?{2�s�jp�	^��ۿ�f�\"`����v�ׇJ��#2z���w|����7V��2o�e�N�F����uE+��\��I��5��< r�_�/��c�"��Mp� �a%��L���OA~�
?Ҁ��FHR##7�J+*�̼����WN����6̎�0D���Ō����n6������Ebk׮<�)��D,�+n4.������%b{��������7�Lkm���?WG���nlc����P�= ߓo��W�9U�z��ޜҦZ{�b��^�O�P��C���_�H(�\����;���86�bٵA�t�r�n�;��cy��&�cbQ���@����G�y���N��7�IV�>Y�-����� H�"����$x�H�Ȁ�<�ˋ�	E•�X��E��8��໊�՘8౾�D���y7{N�o���&�tr��	�J���ڝY z��I�-#��3�(-��H��?&��<,�h��M���{N3viې̪\���h%sm*;�����)�浈1+;��*Bm�B�r��u ��k{�zd�V���ނ2��1\M �ੲ���cU����g��������c��2�C41W�N���,���O5�y���4���U��2+�'��A�	$ۺ��<��]���b������'w��7,��m�|����6
a���tcn20CD�N_G��W(�
-���i6���2]�	?;� �wt��v�W�2�Ur#��R���e�h�?��L-*��D*��D�z]a|d�k��J/uh>e�E�0t$����Q��g��8��]���iN,3�,� -�a*.�%��ߌy`{u[��l��dcv��˷|�����rr���P)��1����w)��
�t�_�1g�H4�5��(�4�H�Z�1�n*Q$�`���d��ԉ͐�RKϋ��n!�B�O+�ouB���n�0��~˸���]���3��,Ƿ��<����S�G�܇y@m�#1e��䥽��4��Xv2����E���}6\��|���6��Sx3^n���mS�p���ta�K�1�^��?[Y���A�s�Y��Bu:XT*�}��|`^N��+��q(l���+.�m���q���IKH�c!1���,�7�u��������h+��)~��3����	{}Y�{K����ԇ��@��F��y21����H�Eϳ�Z�ִ���ca$�kFH���}@�� 
��@�~�i�v��uK�d�"���
�q1E�V^3���O3Z�}��Tq�1	Y�K��N���L��xèT�X��'kmnKu��A��4�Xv^��^�-M�U\(����c��N�A}�r�2�Gq�*8���|�����nD�*��y��P�:�~�|����_��g��4�B��L�Nͤ���|y`l%2Ă['�}�a�aWЉ@��v���@ś��sj0P�nm.���t�ݹ�?m��$�&_p�؞��)����p�(_���	�l]� �L��)�����	-��Q�\��������@�����(aґ-��M�kD(�H?c�+�Kn-#�1���'�o�xbmIT�py�T��c�27	���9�.�x���,�0��7f�_��p@�H�~��{�P�$�.�^c�)�wۨ]0Q�����x��p�<}��J`�<�����߃�������T��VӬ��j�[�,�<��#.�PRF˹�g��}�@bƊT��)+�Ĺws;�g��'e;���ԙ�~�ΡT�<ӌ��- /�>�o~>���+xW��s܋��A�8�WT77* O�!$�'�X]�Ձ̕h����\=P�lZ���ZX����ON�AM���V[�^s��lP��3�r�)���`��ma�J��`M����%Q�o��߆�eqف5�~�D�ӆ��2�������|��\�t��7n����򳦚��\���]r�5�CB�WF�5`�w�D8��'K,������� ؖ�u��@�N�-�-���H#/���'�&O�L�?��g_A�`!�ѯd���#�V5��SwXQ��B�"��E��ͤ����SV�Ռ���0[�$�}���z�0yK�ޕ�^"�X���]���4?�m����<�OX3��.�v��yڑ1��q�3W����{7�G>F�Vg
	W�YVM�~�5�H�I�R�(ھ��w�P׺���/ݭ�[Lk��_��P	�Vꩿ��0I)�@:�(B�1`pgL1%���]ze�/���+�lJE ;���W��m$�zyb�"�c�t���I?=�$Ok��,�=�	H�����Q�e���!!�9�j��_KFKua�PC�v5��6l܇��emԉ\?����k�N��mIď���(�`���/C��V�=�wv6�#Z	6�K�q���i����@�-�rw��D*�����?r���h.��_e;K�hl+"�� �9s�����)|k���o�8�mu,(�Jh�K9㻖x��W��G;'(W��]��W=3�ō,+�
ʉ����4� ��Ԉ�{��ܨaHh�{#������lk?��J{��h1��\�d~0�u��6r�{�L��ѼvE��Uú�rN���n��55����]:û~�h
 ��¥�Yw����Zĭ�E�s���CZ�q�oe=�w����$���O�>9�鍫�E�5d�Ůc]��2��&&��Y�*�E����qj#������i�fbua`������G�e���M�{Rܾ���"��-�E
7��n/jl�w���VȋD�������������O�Z�0�/�� �fv�޶RHͰ�ԃ����RGh���U�7ګ�p}�I������T9,D,q�P�5��$�����=Ѱ�px����W����Tw�Ȝ�^j�W�F̭�k�k��y|�vzs�[��V��o�Aɓ�:�GB�{֔�è_ǰh�ߐӌ����.���L���ʳ�Z����B���jR%U%�`>�T�t)x]�<������{�1**�a���f��Ur ���(����	�f�R3�F}�8�gф�O�����b�edj�+��C=z�N�O2���Y� ���ĄOǢ ?ez[��Z��Μ.��
&�ʬ'S��Y"�X��GD�)���9�S���vXn���ڂ�����O��"�l�� r��~�(���4!�����'�op�����A������/��쑵��u�Рx���s|Kh�ȡ�W{QoF�F���'[���������b��z_ߊ=��oZ��Z$����^X�f���m7P�p�t�Ĥ�UoC��Qo||<}�P�s'D̛����
�>Y��L�X�7�^�d��kU�3���x��'�1ٰ[�a����i�
��̯'�P?}Xiq��\y�\<��=䁕�e<�}a>RqKD���n��MM�����b�w��AY돫��^,�+mq�fX
�b�B`�^�x����(���O=��I�J��_�@b�����?�~o���l��<?�������dS5���,�>1� �:�P��'��)����������+.��ǂ&�{�� ����>dǣ�8�1[w����N��l_�$���5KG�����p���4����N_�M� e8ًX��������9v�ե3�˫�,���	C�L���=zUͧ]uʀ�L�a���'��=�g)�˙��2��2��ԉ��ŗ��	6�^�� B�iٸ�k���3��%��[}��	<���bC�z���{�"6�]����grd�T*������X
�iW�u���b��c�" u���v
�-SR�i`�l�����;�y�#ٮ���'W�)�P��~����6Θ��)� ��-�A��r`�UI⊨�Xв�.��(�ʬ����?`���1n����}��G��+�C:�p�ǠI��~
�2�w��O�C���X���8gw�zo^�e�Y���7e���!��T�Xl�zd=��kL�D��?F��' Ȣ�@�lG�%m��m��UȂ��Lu�|�aĝ��V�+9�y��%џ�*�tM5i��n�Uk�Zf�ҩ�걂y�be7��# �9�� �F�j���	�a4F��\���1ī�=?Y�E{��.I���X�~��x\I ;E�p]�s��ˬ�=X%��e6Yހy4l�u�5���k6�MzM���ZM�S�kZ�G��)��9������3
��G4���G�|R1}��+��i�x:�����U�0��˽�z���9)</�IM�`E-�X��WdR@�^�i�na4� �w�����3��]ު��3��l^Z[}��ZR0�pk�h(����/ÞF_����V����Z,�:�3�;�b��6:ߕ����v"�sy�B����z�\Ϯ���2�F��J@e�. ���@r�����̕R�B|y�!� qu0ws����(sR���%�{��co-!�0����oT!b=B򷳝J��'��l���⺍9����z�f�JL�ceN�������J|�"�1-?f���P�I�Ye,�����ϞçHX{_r�ځ���"���R8���U���x��d.���P�b'g7 rǝ�D�,����V�bpHJ��!*fC�-���c�h�)1*�"�0�a���G6��(�1 ���lx��h���>M����ωhN�l��{츑�y�
���u��^��4wL<;�NeFs���m]#ۘ���O�nq�l�k!Q���'(�'����������}?��d\�W�K�"��1S�
U
$�|�X�)3��%�`~:��un%�QCeޜC3@�H�
��b�n�fV��r��&����ֽ@_>Vi��R��m^���j����+֌����P��l�;�°�͟�ũ��~��ٸI�pE�{<���@�v��耵��7.g��d�Uٯ��ߪ�H�B��Qn��1����v�T����?Ku��(���g1E��S����x�i���Q"��I�=?K_dK�w��\;�I��T�(��mH�^W$�+�ط�}6��\㷉8:ʏ�2#�.��m��mN�e�7?������5� ��e=�e}'�z�r�d����ҵ}Q��_7:����'J���ߔ��.z˴��9�ڃ�"r�
�ڬQ;����Š��C�F�,�f���4�ڪJA@����hT�C��*h�]""n�E:'r������H]�g����P	+J��Ixnq�m��;n�k,ɸB�l�ڃ����O���[�$0r���by6�ܪ�'�ݨ�Tq�u���������_�!�$ؼ0�7�Wx��.o�Ӓշi��V��K��eF�F_G��n���(?�A&�Z�Q2 *`�f�@�lN�Pe����n0}ߟ2k�G��g��!�UP�!Mƌw�7=�{`gi�͡=�D���à��q0 ��:#����_��8U!Y�&�h�Ilf1Q3�d���sN��� ҵ񤉽���g|Mi7P���	�kv$fr|*���͛�Tʿ�;��
)���|8�R�����vBB���a(�O�Q����B[��0}�(\1n��ʾ�O�'h��G18�L���D񊱘_������ �e�ٗ���Yq7�;�'�b�Q�@��*]�cP�9�Ku����0T���
7�:����7p��X��9G��ղ�w)y�w�+1x�^[k��JF;��yB�]}����ˤ���܈�H�/�]�����o޸a�{�Fp��\^��r2��1��E0��ˑU��9Ju�y�/$����iҚ4���3�+QGNl\�cԭ���c�o^��La���� Vy����]9�tl��y.��e�Om]�[�&�#��Oh ��@[2��b�RԠ�A�ȵd�v��`��7ڿgD�����c̘�\�/"5��*^%�I,���J ��7��7${��&��"�uY�3'3f�Ҏ�lx�M��_'B8!���cN���x�ȀL|�>��X�p"�C]kZ��\>�����;����#0���̍i��R���5L;�J�W���+
 ���1�ï+���F�P��\;��V]�7��a��8��]1�\q8�u��vy&���������`��bG�`T��0Jic�s���)��pе���� �}��r��`�^%��ur*>��� ��A�Zi,ƍy�Q����CN�L���:��j���v�-��[}3{ǋ��]#�}V��+C��/1�f�8�f��� Ed�T�´�W�k'pBL�'I+_K1��[}�k�F&������ہrOȩ�?�����g�j�m\�4�l��$QӊN�4_�b&�3��p(n�f�o4H���dg?G�"������KK����p�kf��ѳ���D<]c�$�[�h>D �"�$�����J��g!�֞l�?��h��j\��O�Tig37��3�ӿ4.����4���D� �s(��q�l+�(}P` zmi�����lg,yǡ��Z��a�%z�6}��8ZH���'@F�7ٱK��:��H� 	�fyG�)W ��EcȢ�|~z��O�\��/On�	-Ϡ�`4��9.ꛦ|�T�����:d�e�E�[���BӤ8��(��)O� o��
�$�)-�3�l}�4�Z�6�0��hV�W}���B+��{���#.�#��@'DΤ�ȶdV#y�0s���C��M�:��'�Mwl����Zz�ڍg�dDt�~5H��V����І�=kJƻ[<�ճ�#��;��T�˗c/hr�V����/�OZ'�28�lp^Ǌ�c1��Q@�ٔ�4:^+�g�
b\��!�DSH�bd\��Y�KL�Ӟ����5S��b�ָ���R��G��o*E1p���z��2@kx\k\�2�1l���bY������hG0�2!?�X� &��H�Q������!�8l^<T�F�)o� ��FŎ̢�7ݗ�JtKmQ'h��J���|�o���R�!�P6E�H��g&;�wJٖD�+3�r��pj��b�OF����CI����d{w�Ғ��y�����Ǔ��C�����`��1�j6�1$�/�v)\�lx�A���	�+ `ݻ�����gU��������8���Z�h����Ӆ�{�S1�e�w���?��4d<w~j�a����x���Ѱ�_-8����Z!�4�,&�{�MM/Ҹ��%� .�&*�"�Xf�5�}��1q��"��'�2g���1�жB	Ĩ.h`��rvqCd9�u��0�E=j̻��(#�"~��R�I��2���+I��o#;�� ��������q��Hʹ�b߶2��2P���g��e!T�@����!��wA�d��r�\/Bk/�]���RՅ�nd?o9B/Qn�1r�v�Ch���t��o�0s7�K�*��J���X�kxڸ�>��mbs4�EdA��� ���ި޵��9�>`;e}|lV�F�� b=�|o�H <^�8XC�55z!�����҇���|�����3� J܄��C�}|:����2��iI�A51/���i*�y:�<S��t ���7����!\���b���۝O�y��?:��,��K��L�v}�1�XaɤZJr�z.�"g�t�9
M��5�Ao��uH'�����������������z"�sx�!UNІ�r@�eӕ��4�-&� ��`���O$Qô����T2�v�>!Ŀ��^[Y �PRwzO�Y��$�E���c�+��(���n#�g���� .�1.ׇ�`��>��6� �\b/��I	��I��[]�v�"�g�-X��X,�=���zP�����]�S������bI�e�s6��E�WLq�|����T�!ڒ�֮=�TƧ[鄁�'sg~�O���୛	�8$�O��?[X6Q݊,#��'q+�G�?�������@ȶ�z�:{#[�[;��ˑ{�'����ڗx��7������I�~���@��|C��B{�>�vgR�`��;�W����A�!K_v� 3�?���97p%wsh�ku3�Ǌ*�����
��
�0���;�[���k����M{:O 0�|���h�˱\6��#e�ɋ�B�Y����t�oo��u��m����_�OX�of)���{�>3!��b�m���Vϕb���Ļ0�4��P�^��L�"!.)�;��#5n��K�������Ew4;3|)��]DW
��L'�}DJ�) !����It�4�]��ބT��OHU�b��y۶K<���5כ������T���C�G�D�(ʦ�DO�9���0���o�5�~�(��11��PR䛽���W�l��6eu	+fm�7���o�0�l���Bq���#�l0�]L��N�1���y��rut7%Y�k���i�??��W'm���L=�� "�򬚆���Xbp�u�!�����qq�p۠�&�Sn� Dq�sHyK��_�"Ҝs�n��<�ɫ�>}����q޾ޓeL����Y��J,x����G����dRj�X]gE:P�t�R *_}� �>��Y��7�9��/���~º{�UHk�<�Kf}�w��)q�����w��0�Ϭ���Q�ʛӌ�=�i��x���W���_?��u�����7�QD}�bg1��b��P�����ʵP������\p�Y?,.]Ӌ������;�6���p��	�a���(��j��k���r(S�>x;��+&�v�A]�z�=<�����4# ����H_��K��T�e~~^����A_�>^����ԂO���I����P��#T�������$������k�GâtRܤ�!�ԧy�� 1���x��I���c�2-b�iD�O����< 1�sE���6-�má'��r]g{����l~�F�曈&��!�Q�C[�k�����y6� ����o��wW$&`��xj�qH�w�D
�ٵ�N�?`���]s�;S��5^LON�S�Y��.d�ds�9����p���tf��r�3�Z�_�ܩ��4�(*FQ�����4+�:�a&�5q�T�
G�����~��֩Z9#v��������Nm@�& o�7��дC�aAEn('�n�,uu���!k�b	C��1G�;]�E�	(����C!������g"�R}�<-���7���:��흤���,��_�L���j�2�O֒bl1M����TD�6��\y^&Z*c�xs�j���{���R�k�=\m�9��jZ�b���&�ooJ�!�=��'�^���q�,�����2�)#�?y.�.)%�6*W��-'	ǐ�$P{���>�Mi�K~�)�EEx��#��R��t=���eT B/�p	�-@s��D�u�?�3e��Z�|�l��%w�NDA�qI�Z�܆��JH�X�ޒD�I��*�",�������5�o��UPSx1%|ʕ�*�~��	�'�zZ
?���O�5�[����Y���X���0�%�@�:�d9+�q���ŭM@d6O�����"ϖ�='먤vK0B�����]�N�iUj����v���`o�#Y<q����Z4���)�RFC�@4��?��,�mX.z���J���T� `��/ź�F�Z���w;�T�E¥���X�є��UL}D	s��dE��B����L�:ʰ��O�ꣅ��#��.g	P��ԤY	KRyy'I^�l��1�P�[�	�x斚�y3�3��c�c	�U�^&���P~�R��>q�K|�B�ﭳ�K��;�)l�C��<" ����g���z�?�;���$B�+EĬ����i9���G���{���G�.6.$���K�@(�c*%Si}]3U���-G�N��ݦ?D<�{��'!h��w��Z���#>����,W�u�:��6�A_�72��B��zO�(jj��q[�|�G|�{���s��#����h���x;��<*���9�%��N�����kS{|���̅2,����u��m@g0�+p�$�~_?��T���������M�1�n�y��KǦ.��Ks|8��~S��U�|ܙ����������[�2�O�B�d��E��YLi6Hó�C\QL��o�|iy�)��1�r�2)��r��s��� �����f\�fjE	�V���Y��G4lq�������5���_l�j���yV��)� #�egġ0���t��6���ؑ���~��s��8	`�g�~�#P w(X�c�"i��8.�[�B�|O�,a�g. zfAx�Ңt�4��}q��S��p�`��~4�D������A��x|��K�t8V�����Ϣ�H��ƚF0w�Y��o��Bǐ�p����W��[��i�,t8,�?�W�AS��]ёA	�.��8�L���"�U*fJ&�U�����}R#ݵ��9�l!N9ԡ%&(��?WR=� ��Ҕ��v
�q��]M�W�Z$�D��� n���Z=�s�6
�/��e�\��c
�� d�
���\s�J�4HB����x�v�ɻN��#q�<�3N�^=T(yE�\�o7��\W�8'؆����nh�}���[[��v��ܢb�Ѝ}`J?$��.�_r<}O���i��p�ftL��eu	St��FЀ��kW;��>E���-O�M���[[��۟Sg�,޳�z-	�P�`�,L��ة$ā�[P^���y��a]%ް��ӄi@w��ƛ�*v�4�-��d�ԯ�Q2�ߨD�gT�L���X�p5�@i�� �X�S�W&�W�B��(���{¼G����`��	֥�{�\况3�p�W�b�&�ݹ�ߵ*���Μc�IB���~~�=�$5�ּ�wX)Xx��#�=��r�����m�ů;f�\�����ߕ!�	J�^�j�;��3�Qa�TM�l<���ń*�f|w#�w�]KW�Tc��f��bɼ>ߢ�@�-���B@@T.��i1/q���@�qM�5y0�蟄W1ߛ��i�}���!g��;h������wWȧm0��L�����p�Q����
���ٯ���=/r�'ŊݕFȫv���@�Ц��2���0dp%2���TR��I������A&��]ۚ��|�Z�!��rȸ �]���?��\�GN�Ѣ�,�����*;=4E��Q��D'hq�Ӣ$g�w4l�R9e&Rz�kE!�ܺ�g!�pb�׫���	����;(IT�?�J������|��d �*	t�Ű��=���Q����~8c�V��Xeɨ\��̃/�U�ޥ�²XZ~�O����!X�ek��4өoo� �f�x4pK��!�O�<�J�>yީm3��^k��R�yt�qrX'���RB�8|z����*�r�*4�����������G�
�+�Ӑ�%�����d�
wT�j��d.�Yޚ�D�����=�� ���*���j�e-�Q�"���HDJ��o��/�	���	�?�`T�zߔ����$���a�1����������&|$���GǮ�8� u>�ԋ�}<�t�ʘ���t
v��7��X��_0�T7��.�[O����o��u��gw��Mq�j*��B$ Mك;{I.������	�1�QP�uZ����وP�s�g
��E_~��,���!���9©g�t�Lg�Ё�\Q22��qiw��i��Ƕ�(��=��I�T0s^�b,��ȹ�#��T����X�2jR0�LJ
i�!F��qu����d�(�Q'�cH�q�@
���O������%\FH�|#���;� /��^��\ʔ,�36d�J1i����ޠ��z!�'�:��Y��~��b��-��'l�	Ry��4��3�#/����?\]l��(ߜ�?ˆ��\țFņNb�A�5s##�,�i�7#���yMl3�x�����<J���n�Y(R��x��KYQB�N)��aJo�D@8׶�B��3C�SzΞ􊭲[QC���DF���c~ ,#����h�1V�b�|�ʒ�7�Y\gL�tvq�a��Q�;?�A��R%_2�I|�lp0g��g���cw/�����̅
hA�B��#_!g����u��5��d�Nݙ5��]���9�	�6X`��TV�Yz��F"����w�K<på�޴^寐��e�'�c�[���b$p�>�ck����|}l�׆z���G���<9B�zé���UH�8`:ݿFJK�K�wRia�0H���X/���A7qn8'����K.��0��J���H"ʯ��C�;�F%͆�+��I�N�agNu_����[�tf��l�+vb:���M��̂���~�M�h��^GN�0���2�w|��9fL��^�1��I���m=ssKV#�[-��,j뭇s����4�RU
0�9�]���{m _d�0��F?�ˤl���,�bJ�OD��i����%��LJ!c��[���[��phB*rs���}�a�B��Ni�98�5��poh���!���z� }���8�C���Rxʅ�
ke��,�������K�9��o�~J��EHi���p�[�@�s4��"�5����p��#	C.��',E��y�8=�-w2��n��̺��?�b!�n��~�k�aN�W� �{�E}TQ��z���!�:)/	�%6ܭ>��H�لױ��#e�R�E$��F׼��XLM�h$z�ꆯ[l�0����0䶻A жP�G���K����RgT���ẹ����+���@˝<a�
��U0���	�ʴ2�ܖ��q�4BG��`��80�Q��$rp��z\L�����!ń[�f�ޝ�0s(<�Gw���w�o7��U�������i����"�C�=�	��ۇ�X!#� ��#�B?�U�}�z�@I��Ҥ��9ڇAn9)�1�����oZm�D��/�'�p<-7� ��5��c�9z�9�bR.B��R9tl�'d&���׃j�U�;"�j0n�l9)�-"�.���(>6��u7��:�g�X�h,�B��-����"����W��pCFi:�J�RϿ���V1^��|1-I��ߔ#���v��ϑ:�X|�8���o��oh!zcD���(�����By-�(٘8�7E���%u��Uf�u�`�|I��/��F[ƍ��5�	Α������<���
�8���fK�qճ�
��
*F�%�ݑ¦̜X�lm�dL1��;�U�H���嗠ըЙ�Z�V�������g���BN:N��k1d���r3�$�ځ�J4���մ� ��!r3��EDk�7�"x�y����)�S(�q�*>�.�Y��~�n	>Լ^��
1��O}�[(��:eʨ�ܱw�M؉)lv�u�EfpT�r��Z��hF�
�E�(T�� �e�i��¿���=�fu/�}"�'����������[��t;�2�G/2 r���/epj���(��\���'�wn+�>�7��\�迻�ݐ/�N��E�/�G?-l&���(qt�����p�pr���TwS���!L|(a�.�Li�l�l���tb���z0���7�iYr�I��0:�/(��Ku�u�ȹ��"C���θ�4�9պ�ٹ�x�"���Gզ"!�TG|u����p��V��D�a_ ���B�|��;'8hvF�N3>nv���_�ft`�>=���X�%{lh��bh�;��r�/�rM-}ގ�JrVj�.����/ v�F ��rZr-#pf^�O�����Ӂ��nChA��ci%��X����(�b�F�0����]��I[�w-�T	�6;d]�L��dp�4!�Om�t���6��[ڡP?D��0�S'd���2�ǐ<��x���b��q���+�86*(��������f�ݵE��\���I����1_�kf�w� �2�l�+w�N��@3�=�g�JnǗ1o��p�C�u��ﴔŅ��ZٔGI��0 >e��n��1N���o>K�U��ȶ������1?�S�$x�Ζr ��z��Έ��U�:O�Š<p�B$�a5GV&A���l��@����K`$�� 8zI�����vhp=Mh���"S�7-�D�Ғ��}��ܽ�J������~}Gċ�s&6��#@�
��F�\�4`{'�@<@��{�i�6IRs�_JPEyvΞW\#��j�%�b�e�9m�������/d��B��>/uY��#�PY��|B��|�*^"�3n�;�{��^��xm����*v��zb�l����.���4���Ϣ���+2x���E�߶��h��r+����!Ǐ�m�xk�/Qo|I�g���;73���d%g+���f�V���&�XbP�%�^(�ꎎ�D�b�F�����@���9�o���k/�c�L\6��C�_
���H|�hu��ùX�ǃ��m�=Y~��0>���gI(lҸ�<_�ц��:>�p]��i�1� p~N\,�qQ6S~��t��P��N5&�z��!m5��ʽ=P�Rt�>>]V�|&9��	�<9��$4U���W}ya	77VyYcQU�o�DK�kx��S�0]*���M�(�&�V`��Oč!B�+.�M�zB��,q||������s��l��*,�fG���5L����ɧՉRǷQ�O�Kě�%sv�E4w���$����Sl�Cw��r�*|�Ⱥ�P4K��N�a��)~�A���b���1��ˏm��`�c�gy�4S��6MY�1i��lG�"��p4�ꒈ�G����I�-��oJ wu�?�D��H�����]����� ���]j���������-�BS~�=	)�H%Ǻ��J��uE�w񋺅����ɽDJ�Z^��]�x�t���$�cA��j�82,�4�mC��K!�bV���¼.���N}!Y;,���Lս�_D�B!��8t:QC,�(^}7����gm�>u'��2 �EfP5�����c0A��B&��S�f�,�P�1��*��W�m�u�i���R3#H��j)+nY�Jq�M��'/��'=Uu��3Tt�
�%�F>��;���vT)+ƣ�r1�}U�n�
�#2En%�W*߯�W~�+M�c��p�A�s�ed�DS"�=�|RP7�F�L����Wh���I��X�;�Z���l�IV�W��
�-L��*Xc����`��-|A�T�>��k�2g�|8��ȡ�����
��I�.���(g&��m�V�i����*|9�������{�/t�D�7����ScL7�>����6ʎ��O�K���Cx�r(��#��h/7>�ɰ [��c��{���'<��WǄ�z��T���>ˢ��5�e�+nٵ��3Piw�a�k�H���B�:�W%��5��&��54Q~`����t��cqH�<
���i�|r��Ų��|�G�;�u�ě����Q��`�hB�w
�k������U��i< \4Iqc�� �S�\;���T�T���FL��:hY��-�c4��k��8��v�th��^wBR�d�����U @wZ��f�VgNs4�� ��jUo��4U�v�*�Pr���w.BJNx�j9��!�8��uy؞�</�T���:4��{����I�qA�0�Wj����,e*lJ��=��ᄇy �����˹C��l����MJ�03Zm��Jo'�D��:4�C�K@b��3��&��)��DH8Ci�I�)��ğ�-������`��a���g ���J	?�Sz�d0&Ԅ�z'�2�=�����k�|���@�}���H�je���"*Gәn��|m�O���5A~�w�ԧ�/?O��f�&�=��O
c���nS��;�%Py���U��kf��3���`�����_aE��O��z��JZ�(��2��n��u���?,�'X�4@�T}��;Q�E��rBC�����q)a1���+���ç5�C�S�f%6r���U�������`2��6�đX��Ax�C����+�B�Ic���_��z���
 a��@ɾ#�U�T�?�h]Oi�\
�2j2ͺ=��ܷ��TpF�n���/�0����F8�&��gdZ�����C�Գ�)q��_e�"�k�~>(0wG�5ʃ~��޳���$3)Os��S�/�k�x}���=�`���q���2��3�d~<��S�F��~{�q#��E�7P��+;@hA������Ѭ^��>"���r������`)�I�T5�W���-Q慐�ĵ��"U�2���^`�k�z������Pmt<[$�mx�狴:��Ę8,Jc��`1.����]ľ���6*�ȼ�Y�Р��Ly��ʬm�4�,fJ,O��;������Q��ضx��"����.�t~IWi�����]\�iԛȐP��0��ycN�?U���%����ճ�Z���uW�m7��r�*�vs��O)/���!�:͏����>��_:m��}��+�)C��Ԏ��!X�xUT�L�>���A�3�4�bX���OU���8%px��5����̿q9x������X����z�>`X&?}�O��#H�ˠ!��B���ߣ	-�?���Ăߞbqu���PȀ��>x������fW獑ۑ�G�"���r����K3��3��b�Z�4a}Iz���
π�@:MǑ�����:��]��'<a�L����縅Yo[�'�υYxqL`z+��6��;������JQ��^�B����L��x�%'��c)�-Ua�S@��� ���$��ak�շ��ݼ^����Ȏm��T+���-�u���E]aw�y�3�R�� ���FܖM��cx6�Y�?)���(��9�d����vd|��:T�Õ��IT�w�6Eu�n����gN�^k���3�����+B�Q���fM����Ӆ�e(t
r��aL �墊%��'chuk�i0M�r�ST����jr�9��c#��F��3����C��c�mi��Y6�9��(��AH�5���f�AWx_痡x?�JO j��+�)B�/�Ds����Kc{Kuv��m߈@�ޅ�R���)��r������Wy���A�4V�8U�҅K� o��,^��A�l<�ښ�h�թW��$�JAʬ��E��G�V�	�ͼy9�#>�	�i2s-ط0M܈ʫ�,������
f� �D]��<\F�m�$2ٗ�~���:T��5���XBZ=�!�a
�}���3; �uhY'�~��T6h��������/�r��;��SG%�ᠩ?��oe�RZiџ�cd��./)��]��r�.�bd:���}������Pu����ۧ���z_��#1�������Z�ѹ ��>L��C���?���s�!�,\�3I��n^��P�K��n�����$SG1\����R	��ը�wΚ۲-|�R}4O0����ӎ�^����L~�f8n�j�bW��1��u�K�ŋ��b�?S�#��0��jqF��	���z��e��~�?���:V/�l�cYK�</²��4m��<T�\�i�<n���?[\t%�J��6@��P���{�u�\)���d���D�>�yfv��M:Z�Gf��۩�i�a(��&�tK+�G�/qo�v��m����c�X�-�-}t��s�P���m,�E0Z�Mt�lY�6�>�O*��S��lr$��W(�E���/v��r�����������MoT�HZr��\>+NJ��>�L�� ^��_��HX*�1mʼ��K-���B��ˌ�
fǌߧg r�)�B'������?��å� �������n4�Q���Գ�yd���db1)���m� �F�7�0�d�Mǋ��ZR?��	��"r�N� ��{��
D����`�l���7��7���c�E�%�<B[���>��~�%ˀy�h�x��kh�ݔN��u��_������"�⩺D�Ar��5�w)�%Z���%��pzp���,��[�8��xz��g�t]1��F���#�s�ѧ�F}0��)���M`�F��
5g}� ��VDu�5z�L
��Zڃx�-\���u� 4�(���g��x(|��k|�� 1����'��)+-L���͋�OF+���D����6sR�<zE���PJƞ����k�A�v15y^���5��S��?��PU���]C�V���߫�	���gd��Mzb�H�Z݇]��V.�7F=D��S�9�D8S{�w;Il�y�j^��f� [D����E.��;��n���N�=m6u|ŀ$Bz��;piB���,Kr�.>�e@u������l�W�c�˳���x�V/QߝXr�<8��qRĽ�£ܡ^� ���%H9��UYŦ�1&�[�� TO<gVmÈc�3�u*d���p�Aw�S�=�t>��J3^	%��zhɳ�h�3ɸ�xB���F�A�$sab<��%է��s�#H̝�>[~�/(`�w<O踼���w�6� �IE�A�M���!W��x�2�p�A�T=��!��9d�� �K��#��h���C�E�u�1���3_Dm��r3X���wN�Xzܨ��VQ�G�mde2w����nʈX�k8J�G��MțI�*���4+����a�'v^}�5�)�**����"e�t����'�"�n�a�c]ew�.��Z I��.�4>�ݿ|I?��D4̑�+����b~F�U���DߐaȖހS�K�gMM�uA��qԷ��'�cFX�>.7/���ۘ��F?s���1���}�u�3��	O��/r^��s>�CŜ��ݦ��64�k����e7
����J6��(��0LW-.��s:/�ۤ�J��ѱ��6�Bwf1��ދ��M��C��	Xӈ��\.�0c	����ߎ;�n>
:Y�$8V�p)B��l����K-I6O���5��:>��=s�f[�dl N�}~�t@�p��)�_��<��m�6���ɯ	>S�����j���,Q�{Z�es�q�=����}a�)m���H�0+��Dj�#Y���r�'J���l�s���y{=��1��o$���H�{}*tD����0�R8gM�.J�Q��B�����d���ȃ+����L��Ig~8�־h�s4�9�7vTz�J���-��<{�쎑�����x�烓�bQ���7��0��g[-o!�!����q�ǃ��y6׻����W�����
Qr�#k����}�=^����nY���kN��&�*��2 �wd��w��;0|Xi�z�5A	��"�Mr�@�&�t�5��B�� ���Ni����5LF�u=@�P���;�,��̽@���Vb~�����RBzXٵ0-���
.���{2Ж��Ԁ�E-��?���g_�!����'�� �`��X����}�璤Jj�0-�iV�R]�`��#/x1�E��������Ї���W��Px���No.H~'������Ě��!_��c���\I��k@���D��J(P�l5�ST[^�s��}��ܶ	z|:V���#ZP��>MZ��\W�+�#N�O��2P���(���x�����������D��mwd�m9�]e���(���L�Վ�-��Q����=�v�?7jRD.0��q��esq�yڵ�����4�����2���0F�a�
�+�On6��4�`-,�E;cm-P<x�g����)'�r�@�Pl���pqIz���X�A��/�BG��
K�?7B#���T�	�
�˓L��ݫ�T�`s
��a̳�K�
�t�����zd�X�>4 ��߽Y�T|c�2�5�۫�uF='���(s�:�2(�t�Z�=��/y"E������L��i�Ӯ�Q61���y��صV�O2��:Q3���Ǫpo����x��7Y-�Q�RO"��!M"	�jS
�tԿD	�7����C�6��U[q��0\3�,yx�|��Qx�.�͢3bN�6�E��H��FN�;뗅���k� Ԛ�%�za=�5�lä��13#IE{���V�7�8�ue,_X��m������ޒj�q�e[u۸��'^�`O�0��0m����J�����^˕A_�K�'�w�g_�K̨�y�~��m�{�':��V�:�;x�UF�E�z�W5��yC��X1t�C'�9��R�nF!wXSwꐾ��*E=�u�*�2b����U?j���Rd�t��b}[S�T��'-�����} К���L2�99��D�Tg����u{/��T�wsm@S0go���P�L��\%��%���w�bF�s�Z������dQ�sG`��Y@�$z}^��P_�E�,cB��c��k�l� ܚLDx��	c��ˉ��:��kB:�t�"\�'#󕁦]��Y�P��릲}��K"�;w Y�)���dV�ޙ�i�v�(2:�����ն��q�� �3=�M���A�Ź~�U���-D&�ݫ~�`���	�։�~t�D0�B�u+^�>f4M����Յ�9ŧS`\���&�F��pM�iO��J���γ�Qz��*bF�)P��۟~8�"���Ȝ������!���D �HGΐ�=0.Q:�2 �.�� ��	h�@���p#ʧ�z�ɫ�H�H0���	�2ߟ���NH#��h,~�������|߂�u��2���A�	c]ٱS8�u��zŪ��)d+
2�@a��*�j�$��k^��h�ٳ�zIe��a��O�l!2ϋd�ʉ�".��;�S<ԧ��.�y�,�Iȯ�.t�3m��T�r����<�m����
I?J��xC��4o��=-5\���q�_CiSY�s��Ƿ��ɢxO�Fk�R(�H�Nx>��7�S���״���A�"6�w~q�$&���@+�,��ˆ�^��W043����N}׿�My��ڬ��;M����p�.�����$t脋�l����p��c�%"�$�f�3L-$(�杏�]6��p�k�!�z�n����-������0N�Sȳ�� ���*[Vn�� �8����������1b�Sm��X�{�[��F��Mڛ\��#]��)Zܷg�O��)"?n�$���<j`�׹��l���pۑ��	V>�֜�f�ܤ�*�����ҏ"�I�2�� ��ΰ�U'����[��Qu~.�JtU��z�H�tYvd�m!�fk����ć�[񬊙`4�D6: �ai4�\�����ڦ����(S!����f���B��&�hW��O[l٭6?1BP��&�ΐ��jt��B�c����ձ�4o[��Op~_;�iۨ��~�zr�A�V@,\ܷ�ֶc��	��~��$�4��X�i�>dX����	y�wE��2���(���[ء�	�I]jCOrRm��sH\��;%�D~�e��%e�@�L��D�5S��}N(DwSLe�؅H(w�)5�����቟�K�>}j�H��q���E2���=�����S�
Ö�E�*�B�K� yos�*Iٔ�o��{| �O�����7�!ٞQ]fN"K�;I9�C��^!"��M2�c;\���	O=�E�%��p]��-�{ď��X��^�=n�7���E�k�t���-�NP�p����bڨ��]oS�B��2�x�z����M����7S�
2���/ �>(�zG�׌�q>.�g�n�lH��L�B�߼�}�����U�se�_ ���v�į�J \d�5����}�&\��̟%������0�)�Fx��9ȕ��#�|�>*�_Ti��g6Ř�&B�"�'��ж��P�S*�ԙ�����7�ҹ&���*�D�>�'�T0��j��c	��K�s����E�q�vMdx'ү����5חG���tK�A����ã	���P����C�a Dl�Kξ�3��n��`zY=N�A/I j�K}�Y*��#@�\Ɇ��m�{;o�)�N�ޕ��|z����<�y*Vmu9<,
��g�	�-������N�!c���9�zg�8�f�x+p�[a2+_-�|do�ʤ{�^���s������J�;G*ԃ��t!�CR�r�/�mh�J���Ț`&�@=��#Z,SsR��J��4{��V��T�D��RG�Oaa��w[��q$�)�+^U#���r��9ӃغMu��}�Mq|���3]~�U,¼�Hl�~�ϳ�C<=�b��z�8��D�ϛ����[��8Ʃ���OBb�l��[4Ǖ+�hj�1?O�s�g�Oc���ڸݰ�!������ZD%��g�07дwf�:>x�%bS��N8��Zv�M��1���u�b���Ŧ���*G�gp�Ҝ�̋NdIjx�Ό����|�,d���Q,�|��v�֔Ď]��`��SF�ٓ�O���~Lt橕��E(�t�v�t�	+�����ÍEԔ㥐
��"�\��a`00E�t'�M�ɵbc�*}��c��k�����s�F�Z��١���w�ijy�b#�Yq��&���mU�)�n9�pTes�ֽdj�U�K��5��~�Rl{��u���1�1 �|��k����߰�� ~e=�o��癖���OS����J����5S��l��{��7��iϥ��ls8^�����f����R(熴8
�3PJ�\�t�(�fM��f�pR�<{1RG�i�4�Aq�f}����$D�o���8�(J� ݲ(P�[)�a	�Zs�{ŲL�Q������q���Mh�Y�|b��3Y����f�Fc�C����u��2n���`���Eа!��F;��Gc�E����iIZ����-���&9�3�c��=D|�<O*�^���&���DaX��b�8=\�2���z��H��]'	!g�Ah����Ъ�n��!�_P&nb)B9N��$1
�g�n���g�bI�p�g9�I���6�#��7U%���A/����l:w�;��C\������Kfq̢q�K9{��F�؂�̕$����X��ɻ5��H�C�ߨX��o���
���Bg%���H埋`�㰂�~]1���A�;ܛ
D�:������q6 ��#�)����X;�5s脬�>+Y���@gR�N6�'�]�OL�?F���t-0��Rh���S�Hu�������!��y��,�x�A$ͪ����p�I�Ty�$jǍzw}���H!"�����XD��a�y��ZE07	���nw]q��)��0��q���!�P���@��y�&�gb�<�N1�bD��$ˈ<�K���v���m�k"s��炘M���;����3 ,IyH@���_����;A5�p�,�������l'(g��3��!���"����+�>l|���S�Z)H�|9r4�߯��SIb^�׳��:�i��� ��8�@��z��L�NE+�QO�{��{S�>՞5�۰ݨ����|L�q�[�c#�HgA����"�T!.��Xiϧ� a	�N�t�u�����B��V�(���h.�(��Q�B�z7�j�5�-�������fqٚ�]� P�)*�;�Z��YDMitw2��	 C8b�>��ÏD�D��4*�7���j]��toԤ��ɳ���Lr�4���y��r��&���`x? ��A�9ٙr��f�hͿ�B���U�pu���ٙ<å�Vf��RS��n¯4�4��ˑ}V����K�F��{�z-~�Y�?<��\!ko#�i����7�}
7u����+����*SY�N����{>(&�+��^��ݢf��	�Y�F�l�6�j����W@���e��!�ȷ����4CS�f�# n��zS�7��.\��5���7�Ksb5��\�u���g��H0������TŎ��=��_C �)��Jʊ[��9���ԟ�)|%�v�� �ݹw��6��8=�}^�;��D1d�~ ����+e;���\�d��^ ��hs�������Uܻ~V��]�������xgh��>A�������O����\��S�`�|�)����s%��)����P=�����w��E���?*�<�7�Z/�0+�I�]%j*�� �~��2���6XDB���7���䌰֝���m%|�RJ�D<̯n�j\��A�&93�j�.Ȥj+�,4�r����m�N��e�
N��Ur獕�P��R��;F�?��.���.��w������d�`���]�G�3y�:�0��0��?b���M[�|28���⊄#T�9�uQ3l�G�x�g��['^=T��9��E�(C�U�yH�S(-����:�M�d��fSt���pߗ��}�g3:�QU�o�ыtđl�ҧ�ih�;a�*�ͱhmw�g+��"1�A�Z�l��@}��䰎@��+e��ٰ�ڵ�iƝ�ё��33�ۄQ���/=���q��T-��k&Co�\ ���c" ��ew��۽\C�n����[_��p Y��ܰ�����p��g;���m�׋�ϴ��N�!Ҧ��G�N@�9쵌Y�t�G(0��$z<��hWXHzf��o�J�^WapQ��H��y^�Daӝ��n�~���aL��4=�g���#0�;��e>x-"�8$[j}���>�?����J��xo�37�'���W��U|�������:�А��w������j�v��1�k����`$GT\�^d���k�8�D��@��~��C���\�F�K�7�&�'������I����ǿ�k�軜���0���J���z��c�F׫�N�^n2�(�=��.�(��ʒ*RI;>�J�|>#�s�7Վ��H��)~靼{tⷠ�Uwv�g���^��S�Z������|�t���3��M?�L�ߟ�=�P'���ڟi��PҨw��O� I?͙R��]���=��L����>��u�ʋ���U��ヽ,��8*����z����@�����:^�
r��-�-l�F(�UV�`�bFyba�60
�QV
�����Ԕn0&�+�Jh�`��	�-�=�h*���������a��;~�SO[[�M%W��O�]f�U��x�E��Ӿ}� ��^���瓷�:Q>| �{��>$��b�P�LO^�S�����c%�d�@�t����篠�B����*�US��}k���u��B�!!Г���~<}���l���2)����µH�++���C1E#EfE��j�$� Tη&�e��(��T���Rѵ���C�5���& �bI"�rNǱB=|��	�'�z_�Ke�s�dəa����3�e��8�]�������`>��H��Ah�uͮl�M>��Ԗ
O�aK��OGu�w4����(�+�B�)u\| !�� .Ǫ�����S��"t�ʱ����o���l�_�ԐQ@�}f�����f����!��Zh��A�|9����s�һKpG�7G�P���^�s�ӹ�0=��FuƥH�i�u��}����m��D�{�����!~S��y3�i�?T	S��ȅ!�d�wۊ���VkC���>�0N��(:n�÷3�E�1��ǎ� �J��ܗ�q����E�����q
�Փ�_aV9uI!�i�-�V�[z��>��N�D��p�Ș���WG�:�J���0����V�o���B���F3\�
�hh'v|e0�w0*���`Y�ǵ�����R�����>�X����=3�Ƭ\�33��ݴ���.p���0���f�&4�f����}hN��0(?�*�9:u�g�\9�V#t]|:aG}Ce��D�r�h�;-�4��kb� �%��� �������j��,���!���+���;g�o�`;g��L��?�x3�uU������(L��A2��hk�N��?��F��a�w�<($��Nk�{	t<ń��>����Ԁ�l�c��^�29Mz` �A��_tI_ؼ֛xgb��>��,����<�㌉p8�����������e���Րq�����+p�v���=�h�,Qe�;�^��C��������7?�T�<�������O�\UUtޠ��Գ�sc��0� ��2��k>VS:z����UNC݌���|�fP�$">�-��,r*�JqNnhǤ"W�Q�w��R�c����vZ�c���"��6i���YƲ�Qo��Uȅy�2c��RA���Y�c�T)��0�����7Ko�Q�ϼ��,�Ǳd"��Ƀ:N,�}���Z;�Cw��2v|e�ga1�������aaL	�	������8��@���B�@4/r�׍�鑠{_.�j �]Ž?]��,-�uyr�
!�0�/����m�Z2] 2���v�8�F$�9 ���I��ѩ&�=n�	e&�{y�}1�w�Ȥ�݆�9?�����tѤz��P�
��`#��d&���o�M���`�� Ng7#��c�nBf���3�sÌ@�
;g�7��d��J^ ��Z��-+��7�;�w)-O���=/>���k�.	�Ẁj�n^[JLmzʅ���-����>&��E̻�$Q�:�5ŵ�ȳ]�+c>J�� �^kQ�R� b�$,��&O���%�h.�
�&�����.����[�/�Z���A��P͒�{%<8o�`��xYX@�]�\ �ݠ	�-8%OY���FL��]��&54� ��'����j7	WO��q%�wf��~a�#��g@��u�v?�n}�O,��B��}�p4�A�%������	�����<~J����Te��by�,�|�.���#���"��"�0bH��FF�@	�%��rX�}��7�d�����+�;���] +�i"�d]�@R�	�n��W>��mʀ�yԘ*�W�(�s��Օ�$��� �Fϊ't����<���1��T�` ��gi�ܒ���*D=��[�~��gI)H��`� dK0X���R�'�9^����}~�w*L5�� �T���8��P@w� "��V�&V%zԊ���]j��]d���3�.��_?H�$j� ������&"���8:�kP��D43��9��(�E������6zV�=�2�rMld�`���} \e@�	���s���k���$�������q�<l�>;�V�1��W��D��n�_�a��&���������5�����E��@�+i���0�2&䂎C��RXͮXM��|>;�9w�k�{H��E�Q̀�ڋJ�Q�3���2���3F(:�[b=���8��vԜ)�D�D#u�;�����ǖ��b~�Q�F��X�8�I��c<Yh\A#��,�]D$��]r�P���3�IL�v�#\qԏ�2Z=(���������).�� ��Hqy!^{�u{m��Ͳ~�$S��u���Р�߀�Ͼ�.�)L��e3�DQ#u	$(EGɰ�	�a�ٜ�A�b�@�'3mb� ��A�a�;R�������L�����U��4O��Rrzp�tr% �.�ɀ�QO������qX}+$65 O�3/D�RK����]�B���oP��lK�l�uM�[ˣ.:��o|/�ɟi�� �� �x�߶��6��i0BbSHN���|��@O�ʟr{�?ۣy=��!f��z1��֚"���o�ȷ/�"�������:��7��ssx�������8�Fi�W1���v�.�� T)��+Ǣ6������
�((�vA���X����Ǿ5��s� 5M$��:c�61��-/�ʲr]��T�rD�;x�>�z%��&������� B?������#bq��$�q�gA�T:P�}���cе$!k�~
��jOq�Og.��|`�z���^��?<��h_n���$f41$�ˮ'�l��z���"ƈ��D}�����?���C5���/Ezn��ЖABLa!�%/#�G�[�[��b�|1
���o#��X���qG����7�ي���썏���m�[�5�?&�hi�}���XΆԹI��\f{�8����>��f����#J;"/F�UR�|�>\�kS�Qds�# �X���q�p�_�M�q����u�o4��7�|1�s.s��a$i�:��*����FX�k��ѯ��X�i�fB�_w2�K�`Z<�����Aw�˩��ZA���u��)4�l:'���a(tFmQx>^a�
0�t�� ��'v�$�ix�oU�W�!����"�w���q��Ć��`����(�ۊU\��]j�>剏�����#�B�K�K��f
@�Ă��iy`��I�;F������>�P?�)����٭9����jm����\�p��G�
��*��D��U7��6p�9��������3̃ȈF�&#��PG��!r~��|ئ���PT�}��V��Y
��b��T�ŷ_�0>�Է׼�����h��d���V�_+�@�E��_3^���d3lea�M��S�<��z���e8�HT�ԷK��m�藯�A����l���F�����e��w�p��1Ql�fۀ+F����mP�a�i��4c�h��7)��>/ka5hU=7�g�ό�)�����\4�ڂ��[��U�MM�x��_L�61HY9��*�$!:2��&�;2d'��»�����	���%�Y/9���1�P����?'F�p����S>���w�,�wm$/J��x+��T�f|p�>9�/��_����7g$>a�&�9=��R-��8�Y�Z<���Jff����u�\!stVe��G~��&xs�P����A�D��V����WOZ���t�Koh�PT*�e_�ۋ����a�,69F�7�n�eL��6ft����F�����~<ݦ���<T��S�\��c��0�K��;���X��>z����v
��穪rN$錃�HNn�▢�6�Mةd8�W�4
6��'�ߔ7�hK�F({�GΙ�̹ˊ���9�`{�7+8�����3��KՅ�W&Ahi��LPԐ���o��Ic�t����%E�lϝ��n3+�M��U��0�����t
WM�8^x��w��ǒ�N��z0X[҉1)
�e�n������ŸX_�: {���������s�	�y��c� �ʀŘλa�[[�"�������n�u_w���O6�
�9�}�7�F_6׏�P6s��gfNM!���w'�	�tҤ��|^|�;^D�@��i��q����0%�f\��K $��~��שt�Q�Z8�L�${�"Huy�-~�C��RZց;1Z�g*P��"�ʫ�l��I�ʍ�_��,�3wD�ַ����{ 8��}���>�'ݹ�;�0i���N;jSH��_	X�F]-�Ch�z�c7�N�
��4�IO�� 8��y��u�������M��]��v��pM���ɳ�L��Ҍ+�b�S}�����E&�x>`6W���&.�Y�O�Kp.WPC�ƤEK����/�%��'�AL�D�V�X^�����xd3�A�pͅ9���{����s�
Ҁ��r�o� �	Y��:?0��`���dx t˾f^�f�|D���wx��|�	[܃f~��_�eGL�4F�\��6_k"J�&�%�Ô�/����4�L�H�Y���G�X��vFd~H���ŇP�\0OQ=?D�M�f�����W�	(OO>���Fp��}y$:e�*)<�}��K��r��l����s1���m���U��"��N}�Yt����N��a��x�����1;��h�.��?$9�]�Vj����f��}n��Qd'v;$�u��Qs+�Z&Y,Uk߁��n�Ւ�G쿅w�bs��,��A�룏�;P�����p�0��Dz@��������F���;G��(ϳ�����h��v��1jA�tάU�?�^vr)���qr���-���A�h]���2;�.		^űbG\�³Цukr�!��!�Y6a<	nႥ���֬7r,����p�:��q1��ɚ�!�gFL�>.	��� ���z8�0�dLO9N3a��M��^Ʉ��� P��B��Cf��w�8�i?g�6I�]����dw�t��!V=�T�K�Gl}m�u���rj�Zչ�H�S���.8��s0��!U���#"��w\���
z�h$+�YhFhQzed'#(�$ҟ��]��8,e�<�)7Ʋ��d�����o��H`���{)덫]hNl�V��d�C�g*ŕ7��ؿ.,�DB�r� t�
y!	�LogEu�ի������r�H���C���L����^�Sc� �i9�{�zh!���k���+�?=�v9<�*G��3�.�k�7۫�@O\�cV�`�=Il���������/,rx���'3]f��O�Ĉ7�o�ܱE�n�BcO��������s|b�+�>D}��됞]~K�"? ��n���������sJ@�*C���-�>cR�;Dh$���l'�'O� 05�1�8Mx�^�Xn͸_ε3qq��seS쩿��~�q{�}y�r�s���I ��9���;sN��x|�g^���k��S�����!�$'B<����,q�)��_A|N,������_C�G'K�P�┖�	����E��l0��I|Z��{,'���Յ�%���[�Pg�ao��fň�Tn���A��1!�k�y����W	�~��s90i6��Ss�^�|I}8�~@��8����as��@�j�8;�*R}���j�	 �ِ_�tj邜$�?��#��=����!�
�fn��~�&�����yD���&)w\���E�"( y�Lvnc�:h�^G�B�5C�S-��PЖH�x5��2BY]�˄��rY���מ��S�Z���m����ۊ��0�>vXÐ�!�mD�7G�3|���1#�0��ͽ�X���D7
X|�b�t�����W�p9[��j�6��f�@��.��j�˝���+����&\�Cڶ����-���rxW�;%�ӇR]!�b��b�����4��I��
kE�y�*[!���G���6YjOj�H��8��%:�K�W�Vu^Sn)�/�8 \^o��?�mt�]i��D���X?�k1V��{�q�����yO��f�Ƨ>�5��-�1i�Gpy�Z�z�W�t���$���1.�#��|ir�3��o����3��`�x�3B^�;�I|;��l������K�ƪr��}� �%�t���$����qC��Z1h�=0Y{-��f;\���NL�ATs��#;�5�=.	28-�d�Se���d#4~u�h���;�P�P��]|�J;L��k��W%�B荲�ȒK�~T":�%��3&Δv�]�Vɹ����b�&#?��~\��LM(L&�\���?$�ȏ�V釦�bk]]�C8�������ߠ}�cz!	���qȲ�����DL��y��[���H&���x.�/����}Y�r�L-�E%���Qxuf�V�M��bSc;�]�ڎ��\�S�����4���� g�[�h��J��a̅�<�zS
����mCz7ް�vq�<�ņ� +��J⃺��5ߒ\>���Y�egtD�&H�YJ '�A����(mgq�a��D�>���W�R����ŹY����8�#��J�V�3ZE�����	Ye	.K������rU����)�_h	���֠�������:��I��Z#?�R���l�<�_�5߿�6�N�a ���X��ϱ�fs[/��"mgz�j]��q��8�?�m�YT�g�3�l���_�~���ڠ�J)�3m�*�Ԫ���|�&�)[t�g΢O�·�s;:�R��w�\f)�"�0)
��p�����������6��P�}:���� ���;���v�E���"�����T�n;U%h��X�>╏(_�ʈ��c⿦�n����%�=���>wj4�XK����#��7�0�Oi]��7(�,��Zɲ�����a5T��3m���Q��
��rͷ�=]�KN�fU�J�l®���<�Կ�XC(��H6�*�Gn^h�G������Y�l��^Ÿ�.�]bi\�I��#�Z)�>V{���H��J�^��CQ1��r�n�sp��h:����V���^����i3��g�_8�B���h������'����U`� �A�L"��X@��á&XJU�]yAT�'q�BW���C�[z	��-b�VH��ڢ��9�'�nc]>A������%{��b��L�&�!�iR~k�^�%�/�o
��������׀��(UI^ߨ(�㪗�ğ[�v�TL%�-d�1��vG,���J�Չ���^_�=�B�иI��B%���Wh�uJ�0u�v_�c�Ŧʠ���zx<(�Vޢ���׵���W,<�6
���g=�ܩ`�$�I i�4��z�ޠ!����E�z�HM�3ό=�{��34�߾�Հ��^5�2�W�S�ri��rd|���:���/�,2#��+p����b���G3���R}�I�k��]q��xy�;,�����&���0��5�M���jvwS/_�!�SE���Ћg��j�,i�kɛhE�.����l�������cj>yjI8}<u���`*P�xYo;�ܴ
Ù��m�8M��R��3HI.���t�>���Fx��}�T�E�̖,�����@�y�q�^�hB�D_���������3��
ǡO�^e%�-�9�����+BBޟ1�_ID��|&.m�F�����[  �c	/c�)��7�ofR�%�����{'���E>[�׾�fk�bČ�C��2���3h�G�ٟ�||Wʜ"ۚ@ ���������!l�-���6%t�p"���_�f�i]�ӭk�O�"e�ND��J���''U�Q�gՃ�� K��jqo)ݰG�Q~�sC��AN�˝ ����)�t�1#�2��2J������_��/��u�7�kM��h��Ȯ�J�$nˀ��i6ď��˵�狀�2$���Z�Y�=V��o�ˋ�t���[�ݲ�h��3�ߛ��j���!�tv����}���v����l�;�FJ'^�GXvx�a�ev�O�u|Q�D8^�I���TI���D�b��k�>��Ʈ~�z�$]N�@�a;�ŋ�ǆ%J�s|�� 㝝ѭ�:�@y{�]��zP0p���V>=���p��c=���ŭì��Z[J\�:W\Ac��^�X��<&�		J�Ԏ`��0���Vވ��͢B<�ݾme�H�/�Kf��SmF�e�]��
����g��?���f��B#�3���K'�p}z�wt5����sXwT�*��=S�����9��O��/`��S\��<�-��
l4���?�C�CV�If�� �+\��#�y�D)��}?��d�x�V%����B���& v��:*.����;f;��XC�ŬP�R�ܜ�%
���������ʃ��Ԭ{R�)4���γ��
YZo]�R��g��%s�:�� I��@���VNKlG����W�ì,�7��j������n�&�1Z� �-�*�,e$��E�m��R��?����F�/�(�<���|G�����f+�D�{Uqq�6�e9_�%��IY�}R���G�����i+�l�F}�����:��Ƕ8�N3���	&$�����3]�^5'0'�)��hO��u]�y��Z�qZ�[m��6ϡC�y�G��3���&��C��W�����Q9G'��##?	##�沥1օ)�10�S"�o�*�W�ӊ��v�[��P`�F�*�S�
A<>U��⏵Gt�лh���؇m��Z��웱S��.1<h�0��i����]�?'����<�����h��O`
�	�~ؙ�0�DF^^��O�\�w����4�h~�O��������r\ŗm���	���]�zV㮚r����N���(�6�R?�ی�:���w#��]e1T/�i��W�{�@fs�^Ie[I��S��P�[X,b��K��'�*y��*��@7�a��������xA�ì���y���˟.�"�!��P�;�E���h�?��0��G]2�WmĬ�D'�ߊ�!�e��*ϸ�v�xvǔտR�W�r]�T>H߱GG� �>{=��{��9�ʭ*'Qo���\�d �d�y�'2Ng�n,նH؋�Z')��C��a�uTsV�����rl�[�[��%`�l��s�P�1�a��g��(T����6>#ɣ�����
�+c��u߶	�L�n���aF�Ǯ.$y��ft9�"�YI���x@�VP�*����)&� 7�� ���Դ�y���>�gU�:����R�çw�\��_�8�͉^)��r�C�t.eHˢ����Q^M[	���g��gj�x��FW/q:�!u���޽�v����xA2dS}��d��<�/M�.]U�\\���V�)G)~S���!�}:i*qUI|��Kj��/e��&����잶�4=. �'Lͯ�x��+��;{Z����c���7�l}���R�� �pw�$��R��V]v���\$�>)�(��@0+�Fq<��|H՟z�[�W�=��6ab�=�����?qսW}�ߺzxg:���K�q�/Uh5uB ��%p�`V�h�>r����w���>���ӹߧ��SH�_��A뮿5˒��)���v"����k~֖� w����f����=�ŮN�rY�%���lM�O��#�D^#Nc`���E�Qfj���'zI�b��{f��3Чp��'���d�*x'>�}O`\K���VZ >�
m:�����4Id�/��5=C+�=!��n����Y�O�u�0��iy�iid;;�]ś�t�������D�e������z=k0�����¾������ӭ�������\0y1c{.!#0e���{vdÞ|�L�KT[D^���cƴE�i��Z�*�Qލ�CU^��>l�Hf9��+w���p�-�������@��(�� OON�h����u;T�zU�
������%CP�*�����=��\q���>X}��a��{T�D�b�ٻ�{�^~�����Ы3Y9TlF�z	���=w$nc.j���K�7����:փ��Rn���� ˰���/�K+��d>Qc@jj�;ob#���}�q�*];��ý՛�Y�5!���0�>S_�����395�`%؜�=�;~c_R��S)��z�h-Ԡ��n�Pځ�2�T�������j��0FAڜ�_v1�(�omx�mP�B��e&��[���#�pkk����[�a٦ ���Z��j�9K�ڰ�:����hj ����x6���C@���&g�7.�랏Z��GDk��^ �PXb�F�y�G�5�t=�C4bCb�Nk�����]�>�U4#���F����SXʄñ� �ʕ!��.�.�XI-���c�s������G��T�\{���֋���S�#R0�eT�ɐrҐ=.�wZ�J���ё1��8��|��[GՄ���*�#g�ۋ�}��섈��T����~��dQ��^WSl���b�<�;uԐ��W"ʳ���Io����|82�]������I����#��\!��:�) K��d����+�N��J�.���G��շln%�W_π�`|P��_"�n~b�q��o��n�)�Z��_���~m��H�Hy˪��ף�?���S!�$:�qTa��Vu���R�Z#�*��&�u��Ɵ����Hj@���`Z�k=�7�����b-�'��%(�]�@�	��%�6)	y�~.�2.��j������=��6�_7T]`�����q�L!_�m��g���G�%���~G�(�����
c�A�#t.�#͉撟��-3J�#s���/�lxN�t�'�4�)�ZE��㐢尔�3"�ß7�_�Z�[Df*���Y��>��kH�U������{�N�[��sX��I�{� N�
��6V��.��碿���倐����at� ���8$�	��H+������C��Dc?�Y��(���U}
3�ߩ���RhH���z��z�ڴg�->�˔]���#1K!d�O�������m�>];����/����ؓ�	��dx�է�]���O\�6�Z��F�!��)�>Ʈ��4���j�)p�+F�(z�+9;����"t�J�W@� �^\ѱ[�oR�ύ���f��,E��~ct�e7�������ҳ��F~
�*�7�UR�j02������ać\�B��"Ӟ���Ύˉ�F���D��m�̄�W�N�q��H]��EW>���l��;�q��K\i�J��\�;�Ls�Zb�^����X��S��0V�N�ɥID���w%8_��B������	��a�D�����
]�n��bmy��n��z�vD�����Y�� &wå���
��1�'�"i���4ύx6Cq誔 b��"lQ� y��"S�!��x)�b>��;�s��Y<�U�WZ�n���3��\�թ��Z�HЗ���O�2wP��K��O�](za�v0z߀H�Iڰ m��xmWU�Y�
a��-9p"�Z��[�ܶ�mj�t7����*��q����,**0�Z�ju,�d��*����~�*#�ω��"H?X��o� ����%���o�1�n6.��;�kGж�\U���r��i�8Z���dEI[��rN����x�����d%����&�d��=�M�O��y���+���$�r�くc�$�G��O��a|��.o��	d���.#����ur�k�BWpѳ9��%��a�$#?bF���_8���k��:�9WV7c��J��� �n�¹� �����=����:�l�q��5j.��8�R�����#�'ylQ���V���Lp�~�;5�v^ȼ��We��{Ҽ���s���4�-R-.nR_��  �G�okX��؁����aW�θ�Q�s�H�+l�]���vl/����t(�h_B�?�����@�U��dP"��M�EQǎ'8���wQ���5}^���T�6ܞ����V������;5��C�H"ۖ�[_fG�Rۇ��엘>�*D���iX3�I��a�$�g�Ȇ�:�LC��:����a+�|�A�5�y�-�Gu��y��&�wr��c�J	�W�0�>*Ɓ��MGuU;��M���(���(���W|.J�J�a?�s�5B]&j��͡��B��Z����-�������G�����M���	�L"�lb%B��1���i:W�5Ǻ4���X!��$����f{��3:�?9�au�@|W�{Yv˹��y��ɳ���wcM*�Y2�����_`���$�{�>�� ��4�㛷"!�r]�ϥ[����:g�a��O^�:�r;��|��K�t�L$��"��1��;����?��t�9��)�V�"��S@�H�L뾠{��\fE�I���@�s�h��C՝�q�H�'��ID����J.��<����������Y�S�� 8����Z�*�1�zl�i�T����0|3f��T����#/�A�ܫ���������2���X�EW�o�t{���;o�]��Q�J�g�V��S����u�3{�72�(b���O2[�5�h\&�R�Ȃv�p*� n���h+��_����D���\h	T͐v&lˌ%�0��.���b������9��D�H/��}-�,fWտ'����*B�7��C� w����C��*�,2�vB}VZ'�9&V��s��#��O��XB��a<O	�({M��>7ܳ��h���S驀I9S��;#!�$��޳G3����e.!w����+�y|i�O�KBf�e|��Cn'g Z�v*JLU�������*�1�j,��Ԟ��-��9��g����H�RKnNϵ� ���0�k��Q�*��ٌ&��+�R%Ltz��}�!pO�P���]����5���d�����+�C�5,�Y��s?�'kc~�_q��:ύ!�2k%W�B���H���JMH��Cn}p8�n��
	W��V^�$�%L��p�b��u������955�,���#�f�3�!�;���]~"��B�x��h� �-�Mxފ�o��ٸ�˴;��,���_��������A��dH, �� ��CJ��#��n�M,�p�я��w��07*�^KZ\�L?�9�
��\K�6(��N���� Qm H��s���G�S�� �!_A�;�}3S�3��î�+��~���qi<�lK$E=,Q9�b�����e[���
|�M���Zv"��ʓH��[�EW����T;+�E��+P]�c3^��J�4���NB�s����Q(M_`\��6<Nď#W�,:�)nGAh�������b�>5��e�4� �LJ���*��O7@.��	ܚVFc����[%�z{�B�	�łN�n?({�4[f�H�O����o���7`��j�s�����H`�ʈ.�ACIc�I0��#����Y5�<�g�լK[;H��L�@k�r�`l��Ļ]�P̳f��r��xʢ�h ���t��3R���3�Ԭ� �"K��l��#�����r
�\�,����f�@V�^K�`��st��N&�a����h1%�ʑw,�Z�
��-C��"��ib@��rSz�����pg�1b�l~2bV���T��?]�ôևL�A�@�`�A����ڞ����_�!7g�h��!���q] �&|UW�NBZ�9�d�pKg� [_�5P҉�;�Rvo	�>��$zV�]�>����Еb��������J��#�T6L!���Z�x�%ze��rc�^���?�����6z���Pg��<a��k��l.��"��<N�ƃn�X���O฾r�O�E�b(-��cV�m��-~I���]QC!�*۞���*�[���L.�8��)�8>���$	�$�F�j�2���R��b٫鯉���Pդ��)Khx���Jh�,|ϵ�`[��L�[��:�����<���\s���/����h���qj�Q�u�wQ�B^��(�wM���CX����i��[�$֛V���O3��f ���H�������ܵ�%��1�;�I��|ȅ���Ak�6$A~B,w�,��r�%YEQ"��H�n|�X4���[� y��C�ǩi��r�(������R�s�tI�&�ws�qtљl�c��UsFD����k��ʕ]��]���U��`ux��Kdw��Җ�	h��c�}Vr�a��-oQj��I��L���'[	n&n=b��C���W_\�B�[���[Q"�1CZ�B<�<c�^�<0۲7��������z�|N�	�:Y��k0��?�V"W;EP��͡���.�q�\-ݐ�)B��Q:6�%!|W�y�����eJL�����C��;���AW&��J�%	�c1ÈL�<����z�Z����9�Y�Vz��ʖ�W�g�l�e{>�;�%�d�!Uo��[4%Pf.��F�Y�
�H��0���^�`��U��l��Yy�%r���Ed��A1V��WY��Vר���Y�8�Oa�����ځ��S��5pV���T9[���$�����5����Ȥ?�]��i�B(
�kZYB��ܭp�#�zP����� �t��
�3Q(��/�"� e��4�`�O�V=̘s�ᑬ���r������R��9��X��Dp��Ed��������z�d7P#�qg�7�J4�x���F�>^��㙈��c�Hq*�N�e��*��?/�u�2�mY���LrB���;����o`�/���l��A�J=�:3v�C�_�/ߤ"&vY-��<=� M�z��#e%��g!&�#'�K�p�jiP�7�����C�x �}dʋ�(wCx��Ԯ�+�_5��8�Z��$̜��š����FF��Y�d��4�R��T�D��T߰l�̣��fA��p�ڕ�O#�$\�wU��=����+@�!m��q�_�ČD}��'�ҴH�[W�Gr���V�D��QS�"�me�@^D�*I�J�]N_!�UzWV�K\"�x�<��6����[h����Hct��$�|a�\�=�^�{�섂�����.��d�h7X��~���´Z��\�#�:+oV �x�!�o�o�@�ޭs�<�r:��:�/�A�e1'��c	˂7�5�ׅ����|�?��>(^��B�6y����4c��ڹ�N���'��Ir�k��#��x7�?�����Yw��4�63�	�����n�:��K	�ln�-<���@���{B�Uw"��NvP�C�y�4�.{���-`�"`�i��}w�sc�����31������>��&I}GB�js�5e�j��+'�>"�� ��M^ϵ�b�c�_�e�'Οt]Ǫ������
�*�8�G����\��l	�b�ķ�m��=I$Ϋb6�Ȓ"���i�Z-��=�lvF% TC0z��9��d�d�a��L��eG���D
���7����0����]�1�	ÉtԽ"L5�'oZ B�����nC�Y��7Q�.�\��x1� ��*v�v�L�i[��NV'4���Ƅ*3�ܛ�4�Y��X��t��Yt�- ���Cc�ŁJ��5�Z7�"X+���-���0@Lt�D6
yWޚ�_�먁�gLǌ�Ƚѥ��EH�୍�Q��:���9!�2�{n�]���:nf\ue{�K%f6�����^��ݴ��W#Gմa��yu�$s+O*���dP�Ib��O��ʁja��~P��"rr:Y��b2g$ܵ�^f/q�R�j����,)Aڅ�{()���P��D�O�D*H@>��)S�өE����Xm1 F�*z`Vs��}gc. #�<�Y�����-��2/����!��O���/�����	�Ĝ�U& w�*��{�3.�B4����pn�9�c���V���w�L+P�Aё�r�{��,����BF�ʘ�l��(���="v�����Aw�4�]n��]| n���^T�,C��x��)��]���r �&|��;9�����J��H�Y��(rĪ0�X\K���n�zpd�&�ƒYf$���K��k
�V���n���������	Eޗ�)��3#�R>Ȩ�3�t|'��^S���RQJ	�/{���F+0����ɥ*��Co��{��t�t)	��Jzn�i���Y�c�h�;���;�|"9��t����8#�@w)�~��b����:�Ē�\�:d�cu9�P��vn�uI�~��#�Cw�p�ӵf5�-���E��P&����O�pTDz?�rN�>����>����`��Փ.��-׫[hu�����c|i���~���7ԡw�A[Wx2�}4	��"f�%#|D��L4�~��Qdd�7�\�_^g(-աY6}��z*fk~��8�X͓�1U[����E�;Q)��b��+@0���;"��uxH&����h�z&�Ƅ��'p_���U�V��&VҔ�����IR4\�Bw�S��9cE��Fs4�����B���\،����c濚p��z,��S,1�{� � �q�4����j%���E�6[�Kk�-E�yS��-Z�=E�5���#������ZB��,�3�i���T��N؆�h	���v�+�#�;���������>�C �:����\if��\Fp`���Dץ�7]M�n|,i����1s�OL�����X�����5�����k(�B��$
3��d%���^L�{-�)ڎ@+4/j��E���i�:��Ns~$���Nk������e4���a�o��h��I�L�[��m��[�U��Y";^V��ǀ�!�s�S�DS��:Y4m��ݝ��h�'�0]��Ω��G���E����U�� ��nSV�����Z��v�����cPGy֖�F|�L��Q�G�eM�}aa��;��U�r��x��j%��Rc��v��r��a�6�90;!pq�a,����tk���veŐ�b�Å�w`�b�J��&/JEq�h�hi��侩�����s��l�0D�2-�a���ˣ4ƨ�e�mq	l�o��⨺���fob���j��zρ����*[*�?f��f��D� ?~�Þʄ��i�F$���NcXb^^_/�(6O����#�$�DV�u���W��0cXPkN�r�Q�`k��{	����CD��e����/�F]1Hp�0Z�/�F&j�����~��n��xe�z3`%���߮~R��){�������#u/(3�6�g����H����O[��~�	�j�i��0��T赣#e�	�W���#Q�Ř�օg����`Xf�a��4SfV]rv� Ү�e�'C#H�_�;���ʌ
/xZT�+�I�� ? �dvȃXݡ"�@DH �ݼ��0xvV�tB�<T�Y|/C%!XS����V􊯖����8�A�ˣn�jZG��Q�ي�ĭ|��d�Z����L-��_��",���8E��z ��9d��ﮬ܊��]��-��8q��Oe�Gp�L"�FI,yV��ea��rq��B�z����Tۯ�g�g>�v�,db�+���*L�WP�>.yxaB��WQ�2>��}D
�
�7%l��mGRCy�8Y�P&�RI�v49ڶ��ة9�q#��Ƃ#2!���+p�0j�d)I�ǐq���a������ �W������.�:{ �% ��{]KSbw ����Q!��ICf��I��տ?|E�6/��#|LH1߆|�G���4ҟB������x��'&h)����+a�'R� �v��z5#�m6��jw����\vϣ���8]�9S9I�Z!h�a�s�`�@ ��,���� ����N���횏x���`*k��╌�O8���{AƬtfg�X����d�F3�b�o�t>�LSO}?f�p���n=�NJ�����G�:���t!KPrQ����Օ�_<��зL?ڎn'�5��c���:�ؿi|lK�d��/	�ÿ�%戝.3R�����m�k��)i,
y�
������I�){��.�Ïx��Fz��=���&�M�L��J��\�����@���P���ǵdZ&զ�T��Z$�j7���4����1No�`r���>Y�d]ئ���c*���!<"#�̫���f�E*˖����)D#����6Z�3�h�7m���$�����G���z+9a�\#�؝VБ�"{!��c��L��9q$�cX6�B9�����>�������G`+��o|,�S�i�M��xL% �Ē�]�]�eVܑ��z?�����۞ Z���^�j���Y�x�f�|I-}摊�x�^W�o4�U~wTd�s���l�z��6���S��7��!,��=�Ip�-��g��E���e��-�-�����E��	��u`�,��g(A�#����*�WXѰ&O[�䜸�@��`�*W�'苢�oA&�4�X��F���8B��'{j��r���/��6������	ׂ�}������~��vA^�����Ɂ��}ʳ�\pu��_���;��Ld�
(:�cFo��U����c�y�xK�c؍�ߝ���a�XzB?��
O"2+�/�x�zPt��d��ry.����I	J�� }��"TH��[�|���@�Y�'�Qy'L��M���C�T��{�܅�u�vv�����oN�a-�֊��I�;C�j4	����lb@���_#��Wű,���QXu����%lH�������y�ד&2��z+���1e������&<��5��:������Ayh�z��wa��M�`���~�m%��e��� �[��5������/o<������|�Fq|_�e��h��vY֟���L-�ʕDY���W�J��3-������}ݫ�ٛ#���abicz]
*z�K�M#���v�����le\�%�ڬ�� ֶ��;�A,��t����9_T�J)��7ӿ�z @d�g�d�������b�М"K��q�`�8��F�ϊE� ⮤��З�/�x �6���Q��$׾��$�d�;��.]2��^g8~�=�vfeEw]�y�)���0NF�K0�q��v]r�j��_��yb������{,}8���GЇ�;;����gK�[�ӧ�����0��CG?�����{q���%E~���7�����Uo�� kt�j��B�R_��y����b=�'����6�yc1�(Y'����0b����G{_2%z]�%��	����=Yb�3�ˡ����y��-�_�U��p���G&fO�(��8(�� �\��g����Ϟ��zM��W�l~eN�z4�����$8o�n{9Ʒ�=�N��Z�`MMϓ��.�{�u˧�ފ(qKSw@]v����Gp�$	05���k�J>�F�}DE@�N���Ԉ2��1c�.�5���w%�C��I��y}bB�4�����'&L|n�
�"G�1킐:�=HP_N�۷x>T���.O��OϠ,�C��:='�����t��d�~������B��7�N��y���K.|t_�Lⱘq�"��7�j/���5�� ^x�Xl.����-�*tgmx�ȶRSg�����{N�Ә����5n�����l�tS��}?�t�����a@W4�e���`���]�pzd>�4����N9�c�h�$�%Q�g�wn%���)��|h�>�~h@�l@('ԴKV<�)�2z����:�,��S��=��}�)��̠���7�����-�߮�G��N<l�kk���>�4�ٹO
<�)HGN�s��	������U�>�n��~���Z��;���W�>4")߳�k��Mܩ�9�=7�[�����9�8ED�+�|�ԛ=��(��I���*������]o�7:~3q��-���Xu������Dդy� oF^�x�T����͖-N<��S��%䑅=�>jO�r��5\�Eb���Ý�����y����md����JD�wɴ���.C0ԓ�mT�9��-�Z��Y3�[ f�F�3�y��|�s�U�@�h��z��0�q5zƁ���|���ȧaJc���h!.����c��j��jrN(�re�q�4�4{�!��q.���R��[K2u6{�ɂ��Q�0��-�٠
_��ֻ��+��م��VxY�H�����t&��6�i�.^{L�V��*K0��A~���˗�䕂N^da��6��K��0<�ؗ�G*ւH���}.�N>�I��'������%fi�'�1Qzh��@��\���(c��r�a�n���%�2�� �TA��|���p��<ZgG@��ۃ=�2�м�ђ�=�1ϧ�(]��4eo��O�=�Ē��I�Z��qެ�X�#j��r�6��Ie*d2����s�\�
����\��T����!M����^��n�Yy�9��={������T�Dy����Qý�� (�FI��@��99��؉����Q��c�����>��*vM,�v� :y�s��i�+�V�^#�l2@�DOW_#L�U���O�[�v�-�ZW����5��κ�&ݷJP`m�@���ҕ����D�o�l%�ѻ\u�Z�?p�u�v�bj���v%�=ùs����?+�|�b���@���O_��q�p��oV:~pA���M$C"�ð���̵W`���'V����c=g�g��*���N�D���]+�Hz�������U0���.I{`T7���#k�Gᢦl#�G��&�~R�#��7���+"Vպ(\t^��	
,V�ﴄ�O���B.���R9��p[V�4�>��i1��e��i���&dD)��� ���4'G^ ��-!ʍ{���v���"�/9Φy7��o7p�l��편8�GsUo��T�"E01m�߅�w��Un��̴JƸ�2K��N;��e�J@g�B3���ũ|`��z����p`�[e$}+�^G딺Wr.`fP=vޱi�w��1�����߱�q]�b ���Y��F�ma����zLX��m9t��}w�Sx���3��e�@���x�qICu�
l�9���ܲ���%�?�T=O�N;����6�qj����2P�;9�����?'��;m�5��o��z���7qH�������wBjI��^�a�|���¢���	<�RÊp�a�9
��r�J�r�	<n����^��$���<��'O�Ym�F(;�4+W�!���;N���������U�նQ�~�̝�s�H���0�H
tޱx�\b(�rW |����$���l�ֺU�<��M�v{<go�k���3���]1�yy�*��a������%�&w"��ʲ�4�!.@
U����_�j�4�l��Q�L�W�V���6~�B���&q��%�±o]·	(uQv�'8�aT�^$M^��E`::�avDN	��k����k4��ڮ�xxӗ?5RL�'�D�0��"c�5Hel��ω0b�J%�����~a�6?[��q����??��_o*�@�N���3�B��gok���U��������r!������3q}H��ذ�؄v��ڪ������h�� �TI�5k���e�]�f.[6�;�����[�������7B�^]��$�FI:���0�0��ԫ�&<NI��9�� �F�L�^몓�q㪞��'pΦ�� ���������sH�Uɝ�P��*�� 掂�䧢 d_��q��-���\07sE$
���,3�B�����4���#m�fV#ީcf����$�%�𪌀)���6�Z��j��+�Ԝ<T]]��v1~<\*>��C��a�%���i:�]�'PM�h �G����:����$Nm�����*;o�^�{�=?Cs[�w#Hn&�gx��*#+@m��OR�*�nO�5*bN����üJ0��n4�G{)�4�^�˧��dVc��x9�P}����`2i�lL5�B�h+���<�����3|��s$b�l/����Y��Nݝ�ŀ<��t`ɤ�-�:~��&��}�#���ȥ�L���|V�c=�;�%;�,����x'�D03��<�� q�I_�s�Ϙ�na�v��2�wQ��L�l8�,�J�Hx���	�z�,�GHj��=:|��N6V��KCp��Z)m����d�<�>������w�t0��6U�h��v�Hg#�̡����f���X�}����d:�+�H�J�}��J�ԯ�3���C���g���߿�=�
"[[rY	�$UO��P%G�.&�9���F}�a�5S��#2���?R:�x*n�
��k�ޫuY~PW���uQ�db�|���MHj�u�8��X���af���:Ib3���V����E��YN/�8I�.
�&V�2�&����Gn6�!闁��`	�8C��!�#��Ѻ��wwZ��]���_���
�=�USx�tY%@���9l���"��;M�2�Sp�����4�䒇��t�@9���y%�7ɐ�����n���ˁ=�����u�ds`�+��饘V�B7��� �RCGg�R��x�� 1�<��]3!�$���(�R�o
� v�	�5Ed��^���ߣ�5�dv��ćQ���,gH��?�&L�{�n���p����Tw˪:��G�D4MֆI��8OU�Q����� ��	x��y�>��.�c����e����A��5]��RVBT��!���#� ���I9�6/@�0{��?O�k�gx��$���s!	��ߺ�Y�=�V-�}mekп�c�V�% �O2um[H'YS��7�{h� )��Қ���A�L��bi�Le&y�hS!�A���_�iI3���:�װ�.?��1h��LzYOK��^���Ao��I�D:@��4��8u�i���O��$EO2vpc�Wt}e��$�g�-:xA4C�㪑p-:�>�a�p��F��x�8ak-�Qr�����,�4��_�g�;�q�M��;+>�6co��oך�D��r�S��Sa����_�*_PK�����э��k���b��đ����((�R&��\Nq�}S�	�-���f�n������Cc%���:Ҧ?�擿]n�0�f>o�!��˳���N"{���U{�"��Rl�Q+~��f�?�[L�:��}�#��LӏZ�-(C�����)����;��$�8�"�T��ne}>�dV��ꀈ�Kܵ%v�׋��D����Y6��Qg�g�����Q5XV�y�T�:��@�P��Reg���0f3��u�"w�r�oY�<�+�֨��1�W�K�DJ��摮�ְ7�����z�P�l��8֫�T�YY��4h�d�H:�)���	��50�2��_v��\/�x�gT3���89� k�_�X��>��f=j�w�����-�􀎎R�R�3`�^	{�f3pᇅN7'',�$_�����پ��%*��Bۡ*<9նڇ�nd?���a���|�&=E��x���S^�w�:�DDrNVX�sk�HA.�:�ejZj3�~ՏfJSȞ8�΋%�0��>vn�W�4�Vv�D���e�C^l6�B�NM%3+��^��Ց��{f�g4�J8��LZ�!e0�L���Yη��J�ca0"��j����qv�^9�&��t��wO,���B~�]ĬA�E���m%��X�� �-���ߎ�6��}��3�IyAH�'�~\���S�O���J�|��jhe, ���7B�9�6>�kԎċ�c�{6�z0��&��V�Z;�Bѳj�K�߽��v�B��oY>�n���hc#����4D/�������x�=���BZA|�*J�z|]U�O��}s��5>Rn3��he%\���-�RO��>m�Y~V#�|,����Ì��s>qyKL�E�����er�_0W���Y���M\Lm*�$�X��#B"�g
#b$� gR�%�$�1"�r|��6!eT	 ��sA����-Y�f��ThX��#����!{�=f���q�FއWv/ON}M�|,��K�}y�����!�7v���X�7����ު�
8P�zQ��Vr�TTC�׃�MZ��õ��׎��a�|��CZ�^6eqX�R�p���J۴Y�Qņ�2&���H��m(|��X�f]�~7F���#ٓR?��e=��4҆&�<x�RD�5��_�}��M
ᝲ�a�:�X��$Z��n*Ċ��Q��IT���f $3�ۥ��"k�izd��B0l��v�sK�Q!@"��r�צ��Ԋ��*�=���/zc��� yl�1��|+�JP��3G��y���?\\C��zHot�7n���J�{��y���e��`��=���Nc2v����++[���Z��fԴ���'��'_���໚~8�@�a��ǀ��o�P�n�&�9hfuQ�s8x[��j\9��*.\�R�9Vf�k#GAt�؍�IN�]�af���Wk���=���<��І�V���Ik!p�*Έ[`���3�L;Gi��YN �����VO�'�1R����.t���vZp;%z�ʳ�)HIS��u���i~���݁�ƣ�"L��?q2Hv�|Ä2��;vT�7}e��{_|N{�n�j_r)�J��0p���_2�\��E��m�q��7�^�l��ڡ�˧j_�[�$/��^��@q���������	u_A�6��IkQRpi��z�#���by�d�������jND酢��߯�7�DV�T�h��a��2���t�
ᶛ��-�sV������BI?���h�wU�,�*�n�ϲ�'��AV���a�b)3�2@y1-����#t�8��?S*�2�J�F�-}FW�7�g�S�~b-�c �ͷ������yi�\?8rZSp�?�b����i�qBvPዴ[vr�D�s�hĬ�$�/`8�������Ը>��d��]�9���朝PVc��q��Y*&�R���r��.�U+��!���7r!j��\�l����b�������IĤ<�+�F�����gTPM���5խ.�E�ii��
Sii�6�}��Fud�M�+����HQ������:�&{5K��aQI�`j�O�1Sv������ny�����cܷ>���1>�������	�p�!#�p?bq�-����>�s+�������[]�JF-u�,��Ǿ]��=Z
���P]�p5DͤU��2ݝ>�;��k�|9�n$�촍��)��P�H�1�����4��W��%�� f�f���Ԉ>}�B�����z5�۹���
}�t��g�a?�*��,�s;͏�-F�F�}��M�9��_2�C%��n��9�^(kj��s��]n8��ԊCq"�k�Z�P��A�C?�<���V�օ�|�m���
U�7k��;�]��(O!\�B[іԕ٪d��N��74��g4I�x�U������4�X�e��aqI}�ed�
��?�WuSd	��Ȍ�02������� �ڙ|���{�%��7����4��<Lz��h��q������qP'ϝ��b��^Z��Ƅ�Ϧ����x��,�Y�ٽ=���w�����R��ՙ?�9�EDH��#��/��D���*u���Nl�.����:9�BO� T��Y>T��,�$R�&&rz����G��f���3+�|$��=�f1��_�Z�l�Dz�&z�f�����#� ��d�����(~�-�b����P����D���8/���*��^�-�(���<^���5�ׅqg��3Ӵ��D��a4��K8�h�Cr��h��MW�6I�v2�Ӌe2k�z��<Oo��F�8'q�l�=J b����^���Za{'��Y	��
Z	 R*�<{������~��Dd_<7����d�|�T�^��'{x?fQ�ˈ ����u`s.�_��+^
��\3��X[ ��א�+�huk��ÿ#�H���I��?2���E�r�O�$��i��[����v���VQ�Y���Q�p����e�Ad�h��?��3��CZC�J�X���E��у�ɓ�A�!�3� ��#�޴�U��&�/Kr��}���˩n"�������A�����룥5=i#Ib`���	���ġtB��b�_�PH6P�b���#}��tt��ޛ2�*OO�16��Xç޵*�z�m�����
�+?�O:�'1J��A�|�qP6�$�~q�x�����5��޷z<�\*��f� 4�1ݦ����\�� �%�������o��c����~o�m������!EQ�6� r�R|����륀P�ɶH�H[�>�:ѓ�ǆ�$�[,d_ ���!?$߹�,�޿�:R����k�A��\I�~�� l�)А�i�!����NnK�$5��	��ӊ�Y7	�a��~l�)�iQ��&H�@7I@�}����	Բ����.�0!7�6�wb��bŖ�}�����k&�K��v`v�k@Ne���K�xfT}4�U4�]ܹ��5��Z��+��{��U$��4(Q��(2�}g@��B/ښ� ��L0ߨC���z���J�I5�|Ëj�  +ؕ6+�煮`<peV�(�h]�	�Ke���-��B#s�ιd8Js{�K�Dl҄sT��J�}���s�@� v��l�<�B�����7x�[���@�O�%[l�6g&���j���:&6":���Lt��C�W{�PW��l*�-@�����V#��f��r�6��+"���mMw�7*��SE+��/(7/�#?��J�:\�O���AS��k��O@��o������?��gCB��^��U{��M�t �skWf#���l��C!�DB�ơ�d�����݄e2{��>�9F���s�Osw���؄�?�𱀩��.H�C�_0�ϓC�r��h���)��v����n2M|u-1�����A\ =���ԍ�r˂�0�z��'F́<�b|��(��'~���xq4�	'rZh�P]s���Rd���EW�bXP0mt]��{�	73{i�y#9~�B��ʆQ��;��pC���nդ����B��{"e���VI�h?me0�hU6�;��Z�3�U��Z��IF�z�֒�� ?�U�� ^l
mr��G��ӛ �Z�t{+o5͞��38���3N:e�,��?S=s����WJ��aC�M���#�����UK�R�՝ݢRk�mS�����@����M��m*2և���!��aE����dQ�F{�|��"C��~(�Au�/e��`�0���`�'�GGv�
Li�J_y��(\3�E=��*��?�._}3��v�Au�a����#�|�H׾�0�g��m�LF�{�$�2)��iK$���4��>Grd�t���Z���fz���y���<��waD^;���Q)�߼�S�(�S��6�w`��0Q!�o�$C���c؛�	>����Rq�8K��jYX�Sd{ :�V���F����� r�E*Д���r�h?zh��h	J���3�[��#$�rTEҭ�%�(��'8�|
�nm[F��F�G���U�X��SY���טhU �)�X}~f	��e�L�+��v���B�s"��c-QU��P��6p)�$1��ؠ�1F�R�~�"*���l@�.FҠrƭ6�63��ܵI�F�6�_6,ѫ	Vq��~	�s%gK�"�[�[��e�̲W�o���.% H��\��x�7*�gbb�W�͐�]%�c���-`<�d��_�H� ?��"�s�_��_�;�2۴)���u@����}��Kv�xTd�׻X\����E:"p��Bv�� �i��7�@;��R���OW�k��@(���I������u��>�����y2����l�z��������rd�Ғ�z��m�J�na}.k���=��L�ߋ W���۰��aQ&ʹ�@��~8��j����j�G�܀�갋�R�[���5�qě�T�V���J��'���\l.ְ� ������"��}�B��u�A3=]}F�z�L�n�.ф�\�?�T���w:h�+�� ��9_y3;X�4�B�45I�Z�����#$�X;�!�X��{?����9{j�
U2�#�C���[���xw����{�$����:�z!�T���.)�hJ��0���$�˘1���%�K���e�?���	?trF�"��:�T��*�������'��4K�|���q;�Me��M.4��ǻ=w/���P���m�����}3�6>�~4�*���M�?���w$�)d�.���vv"5h��D��j�(ϸ����⪫��o��3�[F��N��"�֚h�:��ʖ�n��ؔ'$����^)z����1�1ۆ���s���ho{):Ȧ��s����lO�\�c=G"�_)�Ͽ*;�n ���T�`H-��0���_���IN�.L���e��Qo
�C�ӥ����=������3+(�����O�E�X3=���&�ꟺ(�� :���{
		F�hl"t��g�zl׆Z|n���P�JN"{|t�:rsB�U��{�X.`�d�b��K����R)�G�q�A7�*q�7r���({��Y���n	�\����y�u�k����o���l)P9�Z������b��$o@n��]��=F���dڻ�I#�{1i�)�_�<�8��h�ܾ&J�'���\+�>5�*��B�g�4��g�D����A<r� �F��4�	� ��e3��>���_JD�8��6��b�=���M�d{eED_9��h��-�4�[[dOx�Yq�i�:�E�p;)�$ Ml�
���%��fi�H8�}Z)	��u��z����ay��F�0{�M��R�"��L�ɒ����0I%?,��tt�F��:��;K�q:5^a�r��A�X�7�\Z�-�	��ܿ��"T�M�o�Y	�g������8�7^�G���\��7�kwD��و��P���$�l}�+�� ����l��wE�NC�����۵�;_Ŕ�j�K��P��lCHw�6R��%A�W��ץt�+.���
�!�q��ά�
 �S��m�5����y���Ah�m�G(�bD+�m@�FP�Q���y�CaY4��+;C8��\^��n�j�~oo�Z�ISlRd>�ΓY���� ��Fk�BS9a�$��<l�%3|H�#�|s���DA[0�3��]ͲJy�Gƀ2�0R"���YI��)��y���5��8f�?+�y��wh��Hj<�	��cy�P{��۝�>x]��I���n��.��qq@�M�M�L�V֊y���Ҵ	e@�D��a��a���h&�V;���(�N5@����/̭������⤇~� �|�Cfq_�>��k=��1��ѩ\+ju���{�G �f�~(wi���I�U7���-���ѰFh�V�7�,,�����'�[#ؙ�B"5���8��l�Cúɵ~e�G_QfE��gF��\J�Ԗ�B��<BX��h�M�)��|"B�.Z�͐ٞł���WŘ(�1-���;�;�Z.}N��}oR[���j*�R8�=�����h�Cf6���ˎ�-f�@�<�{��������`�,sO�Ⅲ ����n���u��m ��ؽ���4d�k�=9l��i+9��$WS�D��2G���$���H��"�9��q�['�K�M�������Þq�s���P-k��3@�{'�p.�asdq�"k���:�^�u�&5��i5f?v�ou�)C����}F��u��hRjaq���K�U��x~���PnGr�2P5�]�;�Sby�_\��K5\�/8�]��@�N���Ȓ"���N�A޽����h��, `u����qvV���JW�Ca�$����h�_�H���_}[!Ts�~>\��z`�x�-T�fO�ynXq��i�cZ9�N�>	�q5@T�w>M�� �)$F���_*,�"Z����,Cc����x��I��o�n��Lדw��"�k?�u��f�u�ql;S����	{�?��xT���=l�ٙ��?D.@���G��"����w�WV�8%糖llyΖ�A���u��mV��P�sM��f\�X����[Qy&{A���]���T� �Z���xr��q�ǌ�!�S���Ri�9|�=;�[)-G�e�Q�C���Z>IkOD���c�c�4��Q��
L�
����i�!�;����7g5a8�,�+�<�cb|��ܸ$���^�G6@�/0s��U���}�E�*�>���%U��K�p����m0\Ѱ���x'��f�ϱ	g��QV�t(1׌ģe�N<�Hú���IL���#p��Р��j^��īmVZ�Q,�Q��A��V�͒mlī�+�������W���pK����sE��rW��u	{1�b239��zW(�a���X�����������L�� Q�&����(oƱK��G�4}Ĉ��2v%&��68~�E۔8{`¤|s���)KAP]=��ZPG@�d�����2Q���ל��C~"� 8�����x���i�+�(,kj�׆�y�~6&Z�G���T���r ��b�W~�PH��-�6)�?�y��,���(�Hx�B+@���U����[�
���s�1d�4@�W�j�+�T|����	/��n��!Mn W�=�SD���Bۍ���ó���k�@9�:��������DEl��F�M_jLY,߲�]m�_ʛe�b�7��Qk!���R�#rd��4��:jj'������%I�C��K��r�&��&��;��o����:FmR(Nä�Q;�(��4IG:4��p��1�Ƣ���C>g=�ՙ%��I&�h[�(���i����C��9?�8W�U��
�;<-�d�?��RЋ���XGg����n'd(�q��dtj$=�l�$wv�)�_~�J3Y9�ӫ�~u���h��J[I�2�;�<=�?�R�_�B���Ҿ���h���L<�Z�.h+s3��=2"�c���O3�qM�PuպJ(�Q~�Wu���sӨ�vN`^t��-%){�JG�8�rɱCW2**��d!���r��{�d��E5�R���s?1~�a�^:��^�'��>�F���Lc��؝�L4׆f_SS�d;b��ք�s�i��Jk8�U�D�2E��� ei�+)&��vl���$�@b�Z͵X�y����)�_,Ԕ�-��/���7F��B#��'7}�}lӑn�ܯA�|h��?���\�X�Ca�kK1
���E΋�F��v"4tPr�PfW�p�'-�H���F|\ ��́׮�������o������X6q~����M�'0
�����{��[�7��o*p��)>j�1� ���P���"_m��N�!E�Pp}h�E~]Ϧ�_����}�,uw�=Q�l,t<μ/9��D�S���ƌ����o�u�%&�2Zo`b����u�*���t�`��w��Oa{1��6�^��x3)�r��j�Fj����Ne����jٮ}��;�<�'v�s�i�J��H�ܯg�����uZ����@ν+p���{�{����T��:*!ۃ=U�����M�l�(�{��P�G��y� �oA«���z����`�\�饈� �����:R�='�])Jv����\-��0�C-B�q\tI��s�7�Ќn��u��c��Q�o��kL:謼�Zk^\|�(��g�$�#����~e�v7���fQ��f�GO�A�O3@Q1�6%7ϖ��Jp4��2	��c�!U
1 �ￜnB��?���B�TR2-%[p'S���a��9fKN��n�02�����g&Y�6���P�e[����EbW��k�a�UHهH��"E����'&�����b� �P�&�gO���^xhq������.	���칿gWQ��FA��H�;R
H��bsJ1%7���YDڄ�[�c�RsnL�0u�#ӽ�&�9�m"8��eR����N���K�q�ϯ
'L͜�[�M2;E
�v�q�vv��ɘ���L���j�~ȶ[ie������ ��6\L���4��1��dQ֦�oP<i�k>̈́= �q̓���x�H�\L.����"�\*Lf{�b�ݚ��-� T\q x��ܑ�Vs^�F�?��g�t{�AE>7>e])��_@�N��^������s������E*K���<b�ƭe��'���h(��d��3"j)���0A�:�7�g�B��[LՓ��*_�Tl=�������bS]�Ppy˲g6�����r^{�~}P�tC���i���ȋe�wLL*�$Eh+	�5�ǂ\.��+���o�2w=���뒘\���nn.<L�����Gӳ(8�99��r��B�t.��D7U�˱�8|�*�a_
r|q�������s\�P0�ʊ�EQ`���S�I�a��C����g�+5�^IG��VY���K�݇�n.�e ԙa{��̾�v����J�r�ȳp�p�����/Ќil���2�����ˍn�@;�l�o����� ��G���͊��un(�y,����/-Ƞ��:�����*>�c�;{�ի�*Z$g�)�5w>���w�J	�d�J�c�U�r,Ă���I��ί����V-���|��&TD���tU��_05���{���J����6A�T��E�R������@��^x�5>?�J|�P�,��7���pM���u����o��#D/�2��t�6��k:�^I�}?�oᱳ�K���y�UG�)�n�V�,���/ԫܾtY��4"b�r� *ۄT�j<�͑g�?0��h����Rڸr��\�Ш�Rz�ԭ_�o�E�3�}$)sr�,��8/Ib��� =%������u����H�Kϛ'��Tr0�(i�L��{�cw�̢%oi�$i�_�f�x�j�|�f����=ҹ!��Q$1!h�'�r=�H�9���ap��j	�C�1|��������щ����Фw�ٟ�q�=ϟ���F������x�Z<h6�橂����۱K�q����j5��7kt�g�2b&4nWHֳ*m��w����n٤�+[�W&%�*j|�濝��j���&�8q\�����<��"q4��5�0�T�EK�$,�����6�H�`v�E�FF�SFo�0}CvQ��<�>v�$�4����ǳ��y(��7�����ͻ��H�)`?d0 1�}`�_�	.u���⮭l�z?;������/�0�Y�'��W+;�*t^ر�9�-�v��R��QtǻBw/��qݾ� J�����kaH?ps6[=� u�˓4�P���K���MN�K�f.���,��Ϙ][��TXW��J��Ӎɔ"1RB��k��Fp�G�(�N� ��D�q$~�@�ZNڬ�Y#3F~�su]�P:�&�m���p9�����`H,Q�����z���+�U��Q����o�wܒ?=�_dqZ�fL�R�S8�Q���|����;�?�;�+++�MJ;����������
��%*���02+�1�&�:��؂��i�j��|L�.��C��y��3@��5�@����J���ٖ��VA]sQ��a �t��3��O�9/��M�I���H�)�<g��$��ѓ�٢�]��˃�m�s��7QG���)��_�6-����-���A���jp�B���[?o��l��k���b�
�ܦ"W��ɣ��/��P&ՓI~PQN8�*���R�brê�-T�%�2S|-�n��֫q��!��.�I��@��2 (T��g{X�H���DIz�S��nW��$Fws���J��,�z���$�˃d���z�FB�2���݁ВJ�bt�n��Q�S�9;�Gw� 1�WT6���k(��3��������R�~�5��A6_��B��S|��.�u#0��7�*��~<Q���d���skEJ��٩BS�HW�.� ���4��V����ORN&G/ �����l�`�:��Yc�R����S xG	���b-c�<��1ch�0n#��b��[R�7]�//4���\�u;��dը����%���(Oy��\S�����oi�0$�v��i�/WkԠ�Ĩ�#
�|��*GҾzq�kN��F&���n�0�v���P7��~�^��k%λֈo���b��ɦ.���1Mv�#I��ŵ��]���Q(�I�[P"
A}�F�bR��Q����������?�ђ�>�����S�����[����ԬQM4��V#/Z��?֔	����c���Kz��y3��v���X-`�ෝK2*.
�;��݉M�n-�5��*���TB���t�쨝�p	�<���)��+ޠ��Z8�/�c'n~�Р�ί�~1��<ԂY�
����A���A�N�V�w�CL�:���}rP/ԙ�u��F��]-� ��G�R.gl�8&��<�p�.=��-�)1���`p�zD.����A��i��/:�GԿ�2t`ͻJ/�5t����Jr��2@l5 �4��W�^����p+��?J�_���VBk$h�f��\��n��c�}q	���0���/}�p�3D�#@QNd~Ϸ2[�E튬Ė���׶�
(�z���.�y(a{�?��1K��=�9	�y#�9�(1T��eE$b�W�B��>7�!X�)��;�*n�M�{ha���΢5�c�J������-�e�o��)˹ĳ��vp��#v�Je$���΂�FfJ�.x������Ƣ����|�� ���0oM�.�`\�	&����	��"����FQ�5w�yD��GK�fJ�a��j�#��-���Պ��G�&c�Ѿ68�JG�����@�6w��%G��~����D+������Å�ZʊÒf�	��f)��2������Zl]��'|�#�o}0��د<��O#����$yP�g�6\�����@H$'Ӛ�4Y�u��߇������ ���dE��|ٝ�������6)C\����{#�T�0b(��>�M	v#`�:���L=�`2��.j��
���U;�|:mr��` ���8�K�[��e:*�?O�]���}3e�������wJ��%�6~��,W��5z���5W>C_���z�m/�[�sr�P��3;?I ��˪��K�����3�Mo�俁��F�N��M7c�M�4����o�Wj�+4S]��ۑ���d�Kt^�\�w�^��rg�a�-I+8 塯ԁP=��F��R`%i�w<˃�u�{6bs�T��x�q�Ԭ�bz_�Z�t������=�n~�$�A�ϴ�ݣ��}�U�ݎ�(��Wd��j&QW�>�ѵ:4�~�q��qH��u��Xu�B�Ǌ*~���L��{�ϭ}gF�v��Տ#h<ڼ��8�@���)1�E���8Nf��\���,��nP ��j���2J���K�u�����(�Hp�f]�M`��)��5,�����v8W��	���$d�Ů)8N{$��J�bi�L�m~�F>�c��M�J(����a�9Rl��7�`�L�w_���ֽ�;�Q�`6\��#�)�ǘ@9Ӡ�\ݛG����qt��R]�^��z$<4��U[���J��� EMN�8�hx��R�$�o��������Vw���Av�:��]#�g�ZDq��1�!�s�q�4\!�,�'F�S=Pa�o�@����˳"�����h��f��o3d�A�A� �	e��d�ԉE�_o{�� 4O$H�9�� ��C��}^'����F(\�u�%@n�^� ��c�6rיL.�	%���-��2p��{ѣ��p����Ē�������C�/Չ�D�x�ם�Ӳ����BBcE��@+ײ`0����NmJj�����l	r��	��/v~ �~7�/A��D�[�2U5<v�W��0�!%��_GS��X8�������m���
�>�~mÍ1������h (��E[������hʴm�OeT��8V}��%��,Hy.̳0���]�0�_��
�է�^|�M=�U�ڴ��0��� �>�+گe��)����������������������j\+~3�a�Yp��4�
&`�zZ�)��耍SK���p���z�.�t��E)�Oվp�M��v ��b"���*���Gm�,r�p�쪲��=Jbp�2�v���k�ae0���q�d�	���E[�$G�R(�d�Q��"�f��k��ԪU��9�uP��}Λ��\��:�M}1���"��H(<3�����0��Tk��]A��v½�8f镙�1l�f��Qm����NW�n�ZđZdh��q��N+�����7�SsY#M��h���Sb��s�/�=��_�J}�*A�������� ��B?L��Wp�$��!�����
���қls���7,hW��.kRU)�h��`�1ˣY�WY��hҏ�k�>'�MYL<;����@�x�v�,41����QF+G���M��DZ�5)Mp3'b�>�n��k�ُ�%6���3�ȑ���! �
� ~��y9��B�+W�������z/[\B����=T-�m�g�>��}z&Z��L�l�F�H���| &3;���Xa���ܿ:@��R���l�2�jEk�|��,^�5<�{�?�c��e�]�	咽%.Q���T��#�o�u��b��a�K�Y��f�����\Q`t(���ZSS
JE�o��-e��+�>!-M�D;@;Xx �ښ�]V�8Z����4�&�0a�]!��"�\[����H�|� � ���@�k%C>s��s���;Q�а��Vs�$og��?�%d��$�����Rv#t�H�[4꫆�"A�2���8�b��U���>\C�Dw�3�%�I9����'��T��F����sK�U�	E���WVY�6�dvɇ��ч��Y[����nFYhO*��&E��������x����޼�y���F�\�2��^w����e��N�іF,�ݍ@>,��NL?���:;�x&�E���8�\y$Ɠ����t���#���Ig`lj޷l4���ZF��L%�� �Ժ��`0`����z���$�5��
㽣���̩��(��@�n7`��y�Ԃ���T�i�4�o�`��������!$x�5��V���W��#ӔQ���ٝ� a]��*MQ9ڃ�U�dm�0�o1��v�i�&��g=�&k4�A>2���[�$1	F���7ެ�'��{՜�k�����P���onJ�F4{CΊ���L�}�H&��"��;��SJ��M��]�w���Y��J��wt��?�1����L�s�%�����tu]��PI�W��6����1tb�#�����g��C(}V�Gw�l��=�|�|�|h�;�3��������<L2��J':-�e�m���}�u ����cn�+��l&��5˻	$�C�S�:��j>���Id�i`8���3���ۘ���d��!�h��f|i�\�U�G��S������)t�ŵWޯK��ߗ�PE��>T�r�MRg�d�;�fHH0����#Kl��{��������I3�!���<um�y�}��ط�%�^T.��wtqt�q���?��͡�M�lw^O#���ŎR��-�]�<�Nt}�qP�v��^����������]��G�G>S����Tڠn�O`3Q]�D�y.�o�Ex �Ԓ����羊i��n��2���f-�"eN�u��:)���y8��v��^\q�ֵ�4������Z?���� ����5���2�v�[#>4�<O�������ꗑ
l}�;<��EK#2�x*�R����AY�&�L��P+R�
�A�U��ّ��Z�,Kv7�ez�:��;�@��ƽ��&����Rm2e���Ҩ8���k���U{5�+�� ;^sY���[޾��z5a��̤���ᄦv;��Ѽ��\W쾈oXELP3T\���P6տ@�W��w��W#�^A	_��TЧ�� ��d&�u~E���:��偺^����01�_ �����vG8	���_ӫކ���ӟ�R�u��� 1�9`��sokXL���'9ᔲ��|>o����sY�%�_# YP�%w�\�>�-i�ZnA�#���&C(�a��j�mW�q�����w�To�H+l�ޫHi"��7��twDýr;T(��M��ݜ]z���}!"%��u"%�,
�b����:�ˊl��"[�m�Q~������Lԩ����mm�!.��G����4t�+��=��⮍�P0���F�  F�(��˼�
R�� �&����F��,�$�-
�0�~�[M*�g?TF�"�}�*Ux,i��+R��	���t�D�Y<|�J��?z=x��:W�p��g���N�`�k��Q#}�	P |���3�&�/	$k�T�}�h��l�s�7��Qv�^$<���3]��VP��ޝ�@)�q+kT\Kb�Hc;�R������:~W�p�eŘd��OI�Ȍ��@���3Ȕf�Q�O�޺`w|��A�id��$=�E��.���^�;u���R 
���o��x��S��->[Cm�Y����g�M�ks3�/o��L�&;�Oԧ��
^�����#�v	�>��� ���U(�b��j�NR�$�hY^n�(�����]���-��� ��W��\b�X7�S*��|G�_ t�j+pD�C)T�&v�+��Јq���H.�<�5t��Y� )F����$�D����q~��a�"�m�@�6�@������T���.�䶲�����.tÍQ~x��=��;�]�5J�K�N鶴K�����r���E~����s�z���#�-��'LMˣ/����ay��3$�ƕ���c��W;P��Z�*���T���b s
��U��U���ڑZxO�󶁋q���s�(���B� ��*ϝ%�O��������w����I�v|����`��@�\-�4�$�����C�]W�*��e�Q�]�z�`��y�oQ���D��7ӡ�!i%����������S)#Ērˮ��¤�����=ؽ �c�[�����r�xq}�>	��Hh���m�H0ȉT{�L&vI`�Y�<��	����:eUrk>�9���M��4���I�gl/ ��Ha=(����r"�q4d��ҪoO�{��B�s0��ѺǇ-r��v�M.�5�F�[.�*y~���,(��A6�(�D��IZ�?�5�7Ɛ�@�����Np�JS��l�S�j<�\�٭���Y�r�5��৑)>��C�^�U�>�lI��ʔ�xR������z�/@=�����Ȁ4ւ�o]ot}C���;6�@e�A�ʜ(0{���<�0��-u����fy��) ](;��l���v���_o���
���\�p9᪘��O��]�?*���Fs�_Y4е��n>5�7���d#�Ί���r��3��at�B������۸K�g[�HV��!\)qaፈAS�c�6e@���������a��&��E<��E���b���>ݤ�l�Ye^w�:����.V���)m�e�A'��,~��#��m�����a� kb��n$
ٓ�ͺ���F�h1��Z�^��6��ׁ� �j��欶��1L�t �)�ià�����Eȫ�ؽ�wo�Yk�� _�o��uw5VF��1��/;�~�ʨI�gS����@M�8�]�O+��kOd����Cs��Պ�ۘ�Q����T/MSDNYU6��'����	N-��X��(�!#�^L��`����>�-ƙpO��b��+�>����!���/��*��	�4i)����dx�Aa�y�^�#f �B�a��g׮n�^~BV�B�8���rv���W' c
�z�t���b���%�U��OX8�Z�!]A��ЛĜ���* ���i��	���?s����߷�K1��{B�1��.r�;R���E,��
i�}���mڌ�\�O1�LF"�m-�+���S�X쿠� f���<��2YYi����C��L'c��^n//��
TR���<�}|��G�4��KL�?� e�%fx�r�0�߻㻩���g�Ad�4��Dʇ|N��(�Fu��j�T���Kć�TO\��@��1�Ec_���y���R��x[�y}ҤV�m�i��h7p'�|�J��s���F�d&�!�`�"�$D0�z/p�TP�:�_���?cP�o��uo�����#ʜn!�U)X��J����4�T�	D����g:Ժ�iw22?I��Iɛ��:�4���g���.�X���K����V����F�h���M�� ������j�� �0d������>�`��"��|��J�l�色.k�}�f.n�T�7�
�`st���L�d�9I��'��C��"�z��|}��B'����9I��:P���"�X`&���P����d�Z����T�C6��	��M��S%_������ށx�TY%W٪<+���-ێY�Tel��U+ aEN���zN�{#vP����H���=·��iw�j���	|�������~��F7�hh;�R�џE�n�b��h�@1H��LT�u�ʌi�� �ޭ��&,�����u8j��2��" wҖ`�XuѮyDv;`W��`�W����5�t~It�\@���1N�h�t?��"��UnA��9��Z~�V��7`|¦q��Cq���$��{-�"�f����sZԯ��k؟q-,9w�"�a��2��ͧ�z���b�/ �iG5I)��(�YU�_�CfI÷Q���S9`<vTL�'���09� =6�r��C{"����a?���qr�k�p�&�~���_!�H�V]�M+��ce�N��W�ha8�l��ĵd�m� �(N�T2Rw��O�;㖱��ڜH��]�L��&�q�oHD��c&]���2)UV]� �o�אx6ѩ���o}��sT�o�|�ۅ��D��r)��>����`pե�mH돇�s�u;C��&��f�BKq\�oE�������O�g����⊽��|�>h��X'?;k��j�������|�S0���o�����HG��B4�!�S+*u�A�2����_4�T7N�ӓ�Ju����R,vG%^`X�6F����Er��it#�EZ��g����S��M���a`8���s8J���s�->����yh��3��ا�h��/��iR��׌e{�� �Z����(����YRZAx�dm
)�v�����"z�Q�M}��S�'$��d6�U��d֞�c0oյF��VK�R��kX���>�Ij΍#�����O�y{E��TSs	�&� ����GabA�[��;��o��蠯hz��	�Ť��:̍.&�4�qa�v(}���V5ԠF�����K�C�l6�^�h\=����v$lÿ��X�0�\ �B�q��O( ����r�1kWٮ�P�n�-v��J
�l�;��x��>ȏ9��U��l4�Q���_~&���&��3�dnZs-�c��G]݌F�9�[2F��s��p؎E�:�X�����Gy�na�W�Ol�P�(���Fx[3�`�|
�@��K�s�{__�-��,Fk�-LF����<��<�uv�۬'i��ߠr��0y��Hj�	bd*�3�$-{bT8A$6��}��/s5rMJ�{��E�����Q�uHxY�Y	��&@w���KQōR�8�-�or���U7��ێ�R7PMI�QB$�$8�҆��ᅿ�F2�E����\��/tt�b�2��H�ش�w��k��3:SֿVr�6b���ʄ���Vs�Er��[<�R�^N����Gô&�<+�Q�]�Ac,����zvtsM)`��W8�Ib���L�;	��vz\Ԫĺ<�l�=�K_Ic�X�-}q�8Š/p�k=��*��G>��t�&���z�]��b�����9�D0��J�;�n?�A>�rh���3m��j����� �@�*�8k�ްJ,�O��y�A��H�]_6��S�S\��yN�i'����bf�1�2��5Q��C��6�������z�����{{���t����E�����;���s�r垿��\cE)�/%�79�f�i���t�Vk��1weQ&R���(EV�%ЬV�?V�['�L-�U���*͎}+[����$�@˂��?W95��Ъd�/�D��e�wa��1U�Ř�YM&��Y7c���7������#D��+��+���4!�g^� �ITf�]�#<dR?�\g�����N|���:��|�FlN�-"�֣��O_l������`�e����Dt�1��dM�\��\F�-7�����9��I�0 �����׶��1W�Q)�>L֒P���լ���#>�%��R�9�UI�'=�?ɂN�1m@�K��\Ѯ@� 1�]Pߗ�:Nc;8�gME��p�5m\�]�ɫ�L��3\j�Q)x�# �-��s��~ND
���ڥì�Q�S�����2)�Ӡ�Z܈��[3���8O'�{���;�Dz᭻���7�>����s�#�
����  _�4y1�̱ĝ{J �>�Y�76�d4U��F5v�Jق�.B�ϊ�nrD�3.9��D����9��Z��CوW��g^�&I�F�� �\��泣�����DE�U��/�6j2'�7.L>8��)�-n��Gρ��>;�
\�6L��i2v��mW���Y6=�Q��rԇ�<������*N����ݸ���~������֚Ю�WJ�X�V�2ZQ�7x���XS����xX�#LsmW�(�9��P�`�P|��U�v�id�������e%��%K"�7�M�s����Nu�7Rg�GV:���r���CTO9"�	�w<'V��O�GL
}2�km�%��ky�����/��#M\����d���_���Q�i���c�;L`�Ց�� �\�Y��A++���d҈�-�(�4;�ء���ό�7
���s���k��Olk��k**��d�-��F$�ͧ�_�u@���nq$�ңs�6�� �v��]���Y����ՋǤ	�-W�8I\zf����9��pz^�L,t
)�V�Ā�����Sm²�:�I4!_��]���w��Z$��>;b����}9�$�ͣ��/a���\:=��cV�a�&��C������ѴDW;[K���!�	����L��{�;P��\Ɨ���s�<l9Ð�x䏬����1�V
�á���N�l~S�Vũ��2K�^`�J܏�YT�]��b JK#����O�1,�iHp[�}����z�����w�e��������Wٯҕ;�N͂�<��:(UٌU�{�����u���h���c"��՚s�C{��ܪD��C%Ӌ��	$&X�%���ܥ1K �$�f'Zx������iө~[mE��7��ӏ��ɧ��ǡ�%?r,�"O�Y�������E=w�'ԋĞvXl7H�l�SCQ8�1�W����2�>�7��L'5��|������9�!8��"49h{��v�E㐳�6�K|��������;P�wG�sr=zI�dBZ����0.�j��1�:
���K Y9�+sv���5&H~1��>�"�)v6`���@����Ҿ�̜�[r|1�
9%�yk I[z�?Z�\����j��>x�xX��_�w���s�ܓ�C��@a`X&�N�Q��f�2��-}�	��	�t�`�y�]�L��+��S8�eR�
	�"6 &"�bЮ-�ߎ$*���5.71^o���4r��bkƝJ��K��'������8��@9A3���A�~��5t��@ǖͩ�E<��@�1�{� Н_�&�#�JhJld "K|�Q���NWY�-@6�q��ɝ:ɻ_lS��Q��B^�Nؙ�|~����m�E�3]�o�K��B\�^t!��jw���=�!��P��4yyJ�:��C)/m[J�:�Dd�ȸk8B��\��M
��%�P$�V�t"����Ǣ"l�E�~�62�R%�QF���]ީ�̒�6A��4>̥2�0���7�p?<�-��S�v�#��	��F���-�Q}-�����uRS�_�o�m�?�7��P�H<ɗ�86��Z4?!&V.^S�r[+�Y�����%���S�y�����W�7O|�/=�e`u�uD[���S�˰p�Tfj�h�C��߱�wovѺ#�0�%�䰆��/�m�hg�>�Ħ���ۉ(���4���AD{L�/������A��:�-�P=��5f��tp�V�}��@V!R�wd�̜���P�'��W��3��>6-\Q�$`�G��l�%��!�����
��e~�8~�f��Or��_�,�����4}���3I��q���c����mV��v���ku�Y�bo�'c�ѫ���̐�߄�TP[P�\�����?�a�؊W�Sp|e`a��K/�T-��1��6R��,�q��@6��y��ɚm�\c�6�rԃ�|������ج�'�t�H�
��@|�0B��ĘƋ̻�c�k����_.@@�'}[^F���s9�KŨ$QZ��r�w�O(sr���C���-І�^v� �Q��a�t�>��&5�ٞ�]l6@O��ҖJ9��dMv�Y@�
[~<l%��UYO�k�U��<�#6��;p���Q)����F�11|��W�*hn�<��4�i)a�n�S�� VdV \�N�sz���[������̗B[��v}Ud�)jF0�D*����U���Q;n�>�Ye�p�D�
��H��g,��W�l��P>�J<��о<t����� {��IK7=KN����� �wm�����a�a:�ݍB+jwQr%�d@R�N�܊�B�?"�RRd��E-���7wA`̨�f�="��H�b��}R��@pιq�'ˤE��ޣ>��89�DW�%����FL�&oO�lR_�'�ވ͠�C��$�˻�'<(�UW7N���aÔa�Y{�S��]֓X� ��"ީ���쀊2��W��)���6��"�S�y2��xÉ.���j�P�����J��x�El��tWazr��n�:��YJ�Vxd�;�,�Y��ɹO�Ox>����A�s�A 5<�1^���]҄�b*�@�Z�K�//�Rh�qߑ;����&�;��kn�R@;A]q̍��U�������;TX��r��jj�
��
;�0k|
��wE�Xу�Q_�i������4!�����Q��%:\�c���G��w@�Mb��8��̜[P�ck��LZO�_K!}м�I���%������H�-X��Ы�2����$����h����yPi��˜�#�X��z8!�����Y�s2Ph^����9�^�����n<��^�~�э��}LO�M~Ru��|
¸���}����Z��[�1h9��[�4-qH�1���-M�%aHNq4��#Z4�::��)��J����kа[C�UO/�)�����G�)��\	���wL����-oE�`��2EP�[Lp��1&�s��|G��s��+G+&�%0�>��`� D`�*
#�0���� ~� �����A#�KJ#�mdh����@��,|de����%?�����wB��#iO#��X.���۹�]�>��q�KMt��/8�E���k�9�Ƃ���N���3w�id�� )���;����P@�{rC��`�߶��2���6���#h�O����t�ſ����/,o#�\f��}`��]2�\fD�2=�E.�����(�@3g��w������x��+��z�$�_�GZ�i{�b��cS�I�ϩh�U_ҡT$�� �`��H�V���A�²��7N=G�UO��g�Z8e���o���8Ta�P���bX�֨�IU%���Ƥ�f�9��˄��C�L���������j<q�@Cx���J����k�Y��Q�oO[j�=�sZ����Q7�!�Y�5�*Xx��X��u��w�'��p���.y �"�����f�XA�4�ygɋ������^��HYw��b�I���\M.D��~�\���@� R���7<�I��X0,��d������Nȶn��\��o��fc�������z��d� �G.pϾI�Y�ɘPˈ����	q�qq�IBy	=N�{mH�iP�7���Ɍ��0h,��=��O
�GШM���v���]���Z<��RF���D}?D�e��rS�[��ι�J<~�n�t�j�LD�!6�q�S�q\h����#vVL6��\���We�)byc�?
ˁg*��z�~��L��!$>ۓ����&r�c���.��m� U��y�
�"sFI�ؤ5U>�"/!Ж�Q��k(ʢ]�(�&*��V�vm���w�TmJ���X������P�����:�څAGB�g��=;H���"��V��MG@j�tj��[}u ��s?�롸�Yc�aq�u�U�K�mA��6g(���n9�H�&c��5��W�՜M����Yn�E��3���)�"����f�*���Sհ5mBi"�!�q�����~���( �#��AY�fE�CJ�|
�h��?�#��Ek~��V�Yi�zx�
J���~2:�Ϗ��.��C큃c�AA��e(��4}1�J�Xh�+����d�1��Eqc7�eʂ�?�Y��r�]�>�vZX/�1.�ݷÎ�^jOg�45��t!���%��e�b�b)���GH:6��]��5����13�����7S���W䍐�����#Z�mk$m� ؆�9�� ��
����=��[����}<Նp|/��ݟ$�(���v���h� d�����F�'<+RR<������+nz�W!�#0`��r��ubu���Ɯ�-�HNrC���(}��UD���7��M�I�����@\���\xjf� ���;4q��[��O�y(��"5�O�f	�+å$BGll���]d�w̙S�ta��?T���Gm��g-��*�ME��9�CP���v>�ue�=W��J��<\�-���R��F�os�M̎j���Eh�okZ�[٠��y��yX�4s���'Pm�ѵ���f�Hw)Pc}��1 $[F�Q�CD�'3c�8#�_�cVI���6���0n�M4#Ж�QD6j��#5��#�k���.P�����T*<�f�ʮMB��&��'e��>�`�ԳUg��ߌo�#�\ʱ�/� $'���<ދ�����軙^Qh%L�C�Ρ�P%��L�9��i(4ޚL��4��]�Xx7O�;�aUN�M����e籋(��㬢�	m����IΏ�&�b��z �&ԡ�U������m�Oe;!ڌ(sʰ:a����yż�j��GY��3R�Xӎ���Tx���6�<�:�s<���l)�� wɱ��a�*�ǔ>��wH훮t���21Rf��c�#E[�IVIRo���؛���_I;�lw�J�*�J�`�
��-�?���~�ϐ4�qy�t)ǺĖ��~>��1�űG�]d��5��
�����$�W���G�6Rh,�k�� Đ����7P:Q����Vyk��c��[��k$i����_G�U�d��@n���	�EG$
���
,,�%M}��tӒĉz��,h[#��@Č��[�/��U�g���m��S�
":����Q���.L�`��KN(�T��œkԡ�P��&��d+�Pث��^��x�1�""����f �`�M�V��H�	��V�H�l���f�	)���w�<{�E_�:"V^�Q%W�wG&ޛ ��� 5r0��{�Y�d�D���~�e��1ݻE4aŦ���S*f>�K�=p(�3��Do��H�V�(���ECH�<fEqN1=���� ����rF�>��N�MY��d�o��Q�����]'g��>:����J4�2?�h.֞����=:��ݮ�^�k7ũo`�i�f�i���7m�Q���6�-�-������՗�Г�G>�+]j*t7�i*S��SX���=�4c��F9D0�Q�H27�C��WC�G�K���Y�y���3S;���zӱ�t��qOXo�ZL.t����W��-+���ZށNh��J��YX�,��W�6Y�pz�0Cu���,mͥ�n����ƮXRs�L���w�����Ԅ�1�� z�`����������T8�R#�W��P�`G�,ʅlab��/gC�=�:���Sޢ��(N�J.�L����H�5�l�D6�1L�#̊/Yb���A��A4G9TJ��ltZ�gJ�{����6����0�<�\]�T���t����ѓr?x�c���ڏZɹ_�_�ԋ�=E��*;aD:���=��������c��E�����Sc,M%�,v@���C�-����yO�)[鮅�B�o�_!Uy��;�<�ݑ�+xȒM���a���r8ed�o���Hh�(��@��� 򃁮�a.'�|��3$�K̀�$lEt�E9隩u����b腡"��
�����s��(M�h�+�KR�g��8��,��k���_���X���da
�`A��}$�O|�%^��̻�����3[YEK�l�jAl��	B�F��ap�Y���3���� �� ��=���Iv{�g���`��[��U2p'�y�wR��uAh6�B�T�$��-�!-S��	���gv�Ӗ��8h���z}����.D�L�ʚ���"_��8��Cw����~9��q�"J��}�-ww�/SCZi�)K�g�z�1����a�F��c	|��Ğ�U��ʞ*%�k�`�.X��sC&���.��?)��
�15[�Zz�ѫm�p{ĽoD\�[�����"��L��EO�:�"gp��,�+V�)ESn��"ˀ+������+��)D����l�Z��s��j��A3���V��-ܦ	]p���h{Pgt�Dbr�B0�O�jw�o�Xݛ���\"m�
I�M�f���L�zu)!�C�P8\�g��]#BR��P��fS�jw(Ѹ�`��z�z෠����qVd�M ������4֝Ж�=�<�l�jr�%A���1�2]�=�Ѵ�4�S2�� �����?�şg����#ӉE��N�I^{�T'�4���ڬQ32I������<�%�	ݳ��VTC	��/�𶛵+�u\���j��^Җ����yI[a�4��N�T�� X�D\ɳ���\b9h�t ��ɁH�>��Jl�`P�HK���՜�?��C#3�i���a�]��,���JC&'����&���";0M��r�1��ɅO�V��@ڪ�xĊ"l:�w	���$@Y)d�kG2܊��c��������[�g���L� �/����J��_��C�Tu1@�N�=0Ɗj��U�x�4A���������q���J��'�S�%p���+s�q>0u�����D
�2��o�
*��;M����X�#��}V=J̌J��&�V;�>�ॱ�[�M#�%eCZ��^�^̋��eb��`KKhm1�pg�!I���D���M0�Əl�HI�ss��Z��1)���SHX'��ϒ�'aH.�'���(�h�;���������;��̜`
��ԯ���)�L"����{�@B�}�Q�]�א����޺㊬�jO&�՞/Y�@	$��Hx#���D�֩O��O&�)p�di�p��G���P�;�/�[/@�1(�UC@y��F&��,��i��@�8߳4�Z�P�F14k�:�+���VN$F9�C(C�ʞ->9�P2s�Q��b/bY�ԅ�5��z�`$0�ԋ�Q�=#fdG�:�SM!���,uȕ����.�Rt�	��`eK#\e��HI2��Q��W_�/��U8�~x��7R��<��}k3m�<G�4��}9��N��h�� ���^o'���V�Sݴ����̌�g0[ЙO6-/Pjt+n�kJ��9���'��ݟ�PMu��`��[8q^0<BEvb�N1Ր��A�*�`�����r[}�[(����Br�i ���+��v%C����Ɨ��چ�l�7�:g����v�����R�$��]�ւ��æl��o�J\u����f:O҆]����=��n����.^�s.0�m�柦7x�U�At2i������mx���P[3�|c>ծ�ڇ�+�M�0X�)b��psCv͆�0����u	G�W_͗�P�p�UE����B@��¿�0m����t��᳐� �ٵ}	L���HK��K�سq^��2���c���Ө�zہԡ��!J�񢾋rҖ>�O� �=1J�������OT/��!�c^0OVV6����U�%�A&�Z��ҿO��i����m]2κ
I"Uni�(ԉ/ R��Vʿ6+_j�K��a[t�e����U���)��^��[�]� ���y#�={Ʀ\�1�}�G]L��X����93ؼ���ur#��U��%.'1����km
�>d$���KF�҂������.dm8��E<�p�N~|u���(0g12Y���	�0�z�ށ��	��|;�.�����R�Wk���"p�r��wZ��^�*R�ͣX!�\���I5x1>h��;n_^��� �{-0�M崕�0m�mw]7DC���N_���r�!$>����.�}˛0�Xc���=�/> ��+�y�I�J�n根�l��+x��#�����V]�߇U�Qɏ�(�AAb�8Kz3�y�Q����v�<p��J����� �b�,�k��>�����^'��{�%�~CJO�p� o$UkbHUv��Yo�Pz�b �L�.��%]�_���m4�ew>�K{����m`��Ȉ�+�s)�f�(m�����GPC�\�
������A�e���={a	P�lYV��z� ��yք���}�R)�?��Ggm�a�*�,�4\�1bA�H>P펤����U8���/�&�!G���1��O^�@M~��g��}Wy�ZH�%��p�bn*�KG���	�0�e���GA��ܑ�hprdq��Ҳ��(t}M�=,�W���^��>-� ���$�1:����< ��G6��b=|7gB�k	h���xD`�y�Y���୶ſ���,����Χ���p��H I�����e6��0��k��;�P��"gy�f��w@#鎘yF-M��ad��9��}��,B�oZd�&���D�
m��qF˅�牘@��VN�G��[��\н���<e���/��,)�����%�� W2�����-D��n1׺�͢R򳨠�ݠ��`��(�Oy��Aco��e ���Zd��QX)��*{W�.?����7�tg*ED�Wt���.�y��&j�fȬ=\�!`e�٣�O��֕����qd� ����TUy�Ldy��H�F�fVI�Z�%i�~��Ǒ�NCg���l��YJ�`'Y!pƪ{2�Ui����E����T��`tV�B�J��-�Q�ψ������VT��+�ZfM���3�NfI�	k`5,Ύ������Y]�@k���/���9�R��.%b4O��\�!R?[(�����h�s������1���=�g��t�:�t,;��5m��T���
?�'�����ȉEBH�3�\i��D�r��5�v�&�A�SA�'�d��J
 �7?��c�����[�~��L��ح�X`'O�3~�f!ْZ��Q��Ȼ�+ri[���g��#��LI9͟7~��g����]#���_�n���W�v�K��3�lOr��4�\o+��R�*y �ݬ�r?Q�n�Z4v��<K��H�O��+4���2��5P�Yum�LQK=�7f!�5R���ͪ�ᆁ�� @��K�Դ����s�R�q7֏2�m4;M*�kJ�����{��mi�v�k��� 7�
L}�F�eZ�~P�Uƍ��O��`�?��@ŅHL�-�L�)��t&�R�+Y��5Hٶ�hm	.�u���̿6֑�*!���X1��]
k�|�`�6��ߖ`V'%2)fA�E�7ǀ~�'�փ��&r{�h�b�ހ#���>�\�=PL�o8�0r-Vq&<�i] 
lAX�{���.{ڶ�Dj�֑KCE&:XR�ol�>�gr�]^3(ȏ/WV�Z�@.e�˻t�Z��!�[	xmXMXV~m�:�3��0mDA�m�1]�qp���y?߮k��57�K�w� �����n>���<E�1�M0#�
�2�8p�*B+� �$4?��)��R�H��4���X�y0P�!�-���"K�]��Q_'uҮ'R}���UY��;OX���h�J9�|��,
6�P�0��fV ^ҠhT<��0P������+^�~2
��$Mu�6n٤aoK����[�j�τ��l%~���G�q�*�X�i,kb��3iY��ˌ�F�M8V��%C��rCX9��-	�8�-�찋�e2ϖ}�h|�Cz�0a�R}�>�,�3Җ{�ԍ�k8�\�U�	7K/�;c�������8+�_�����q��>=m�y�v�id�}q���	b�@��86F�j"V��%I�v�.0
W��j�!��@�X>�ut��3O��?�Ԯ(ه²���p�	��k�����op�b�Dc����^K���ǔ�x��P$
�8W��b&C��iWv`i�{�כ7OAN��iY��R����
YBc鄬�h����i��e�PV�l0�4����*gr2���*�,�!x����|lQ9U�%�	��7F�:���l\��˧�ԛ*�O&�Ho��z}��چ�3rN���0��M�N�<b�E'$�F�?��j3��n�{��$�oF�x��ˊ��wT$0U���w�?��E�B2�=i뼎S�@��8�z�\�>��`,�K�����|iN���E��*
�hL�\��v���H�Iכ`Z`�:V GtzP�� i�⣹�j>x⋤�G����+��������D�r��nUL>*��*m�ν������ү��Yz��2���gZ�F�`���t�Q<F�Z0���p܂*�n3��|@�6�[k�xn�Z��Ə���w����J�:��i��1�oxd������>���jT���yں�;�����b�=R} ��'�Q��P7�	C{����nֹں�F��s:�S1؇�l�˵0>��U�t�Z�tSy���1� v	�֦ u�Ѕ?�<�@�e��F�5G0��˞���[D�v�_�Z�-�hf �� ��ݎ�eĢ�)��c�ƪ�R���p�ìL�58���������vmC�5��U������ɐ�s�(M�$��P��sJy8�ʝ �n�/?�<�
Dn΀ ��I�Kv�Z̟#?�--��OG[Y|c�@�(K�Q�p���������v�M��k���k�x�f�)P�)��}\"�"R���?�@{�17�ӿ����B�z���9g�l���������J������5	�"� �8s�
f�Tɡ���" .��P䖱��RON?�O�m��F)sû\(��l���k��@ ��(c��m�4�N,4��Fd;�v8a��3E�:�������La��" ���<.�b7��s���J[~��4r3מM+�p�r��֘H!v=7z�V+�.}!�*��Qj��4.-0_|K;z�ۤ����a��#�K�������Ŋi�߁�eo-w2o7����!�+��:�� ��t�c�P���X�Y��e홋���v9RJ�� ��bԮm�D?�0�^�Z��8�Q���&��4Q�X���U~��)���C��E���� �LŲ ��:t���D�A����C�Ֆ��E�,Nv}�쭄d��&�P=�inԁ&�+b���\Q�?Q�G�,){�FZ���i����J��:��f���j�J�� X���+a�B0�SW���]�ʧ<F�������@�4W(���-5���>�1��ϑ�M�95k��^���i�_4�T�p��R��j��Q�珞{��v����zN��������J{Ƭ�w�J�	���Zǈ��Kxꧯ�ڧG�~���)��C�~�;H��~F5��d=��Z͐����Ȓ�����6n�z���,��?��z��h�Ĺ���*�4�4ؼ�6Y�PF_�b��;$l���Q��b�����t���ɼ-֯!ԇK!���4g�d�Ҝ�$
�xe��FG�֘U���ZJ�?�Z��~�dg�>���Ӓ�����Řp����'���s*�Sl�5�Vb�~�8h`�Z?w�|ހb���>7��_�ZU,0^`6��ۯN������;�J:�z];�=��rSU�`Lɗj�m�����e$��M#E�>��)����ފ�ƺA����C��Dsѡz,� @��D�4{�:�@���9�N� �2��$�5�9�n�e�s�S��o��k�e�@��M��.L-��W2��.'-$�J[�&^��ܣ�`#����"��=ի��D7��M�<J88)I���2�CE)�dwk�c���sv���MH)���s�0�La���$���Mq��oq��G�~���kP�FKCbd��,z����«(��v0�6[AU�a�@}x��mWvdV����Vߚ=B����&޺^�½>4ӊ�'�-��ۆ�}5�*�(� X��0p�'g���z?u�vbx��������R3"3ٜA����NRxL���%�5-�]f�GO?�*���7⌜��'����Z�4T��"|wSrT����I��z 7��7&��	�Ǩ�a��"mv����ٗ��!��^83g��R�b�m�DܪHu����O��m��5plqЄ�[Y�4�eQ\�AA ��g]�VPZdӢ�Ik���gh����e-��Ǘ"��'����82nr�Fd��o!W�"�{�a�cڏ���"3����D`{��
��S�F���6{~�Kx���ܼGO11�z^e4��o:���a��dy.��?{gm��aZ�!��\u�~UDP�gXE�	$�4��7:M��c[�S�'Ҟ}5r��`c��R�nL��+��ڰ[ޝ�@r�-�1�Q��Y	��`��*�s
!<�:�!S�SL�S
��$��~;�蜅�"Me-x	��c�^䑱�� �!-���l2�$���~�������g���$�ܮ�+Xx��*rj����a��Ql��K������pg�$1��$�6�4�j".n��.,��W������%�n��Ĝ5` ���P^��akO��r�f~��O��`Y@L��m�h�~�g)l]}��o]p�>�G���O�.'�^�(�r��,5��V:��e�'�(��ew�[U.�z��3��xR��k����`�����\�� m�-�U��v[���H���B�;�ѽnD�%��z�V+V�$�tG]���]I�t���l�ɣ�	+��
�H�H߈�)�����͉���}��?���I)��}i�K.f�*�iJ��/vkteA��8-xI�{��I����d,�tS8�$K( �*�zjr��o�J��H�ZA�0�G���m]M&l�y�0fӂ��8^jᄂ8AJ�	�� �}-�zm�����w�x��p���	L���9�����S��LDqZ"�=iH�j�b�����1����y6��0-��ef�d�������Vӧ�Y�ˀs�Ժ�d��͏�I��|�P =k�;�� �>��iX�P��� �r�K-�qM���FP5�_ZT���p�Ae�Q��{'����6�G�-�7@�3��sښ�[2�3B[��e$?�}�-�F�Еd�!!=M͜�P��b�ޙ��S�`��Ƞ����h��!C�����E�H9�&܍� h�+n7�����̶��j�İ��֢�^\l]�Y)$�����Ǜ��6K�㏨���}�aE�d/��^��t$��Y%�+ ۻ\o���dc��ahr��/3x]~�F|�e���|c,�՟0L?O
�؆cG^`�(��	~ח8���9Ǆ&EZ[�v�jE+K��P"����*p9S`�u����6�K�M{�&�s9H%}{�U����b���Z����-u��~�tz���,^�}�p�W�d+��/�u)�|�3�t14�]��q7��㟄�k�\��t��%kd�$a�i�h������\����<��?��}^�;Y|#����LkiS���w��4��R���80��G~�'��$�=�����:^;�Ѩ4�11�c���!�`�n��b	���W�R&�ضW3�]��}�	51���%X���d�٥��#�:\8��=E��e��Pw��j<bͺ�3��}Ը�X�/D��u̊�����`3�2�*q$P�{*���G掫�g�9J��sm3�5�L��[;@�k����`PA��~B�[Z��b�n��Õ��$����]5��Cb��R�5YHE���ơ(��@������y��ӹ�A���s�玘�w@��?vi�-�(�0���_{�M������p�Jo'���!Mp���]V�kR����z��Sd����"�C(ִ9!�kk�F���It*<> X�:����=^�`ٰ�Ay
M��ۊ")Y�M��� ���ɛ'�:�!�؍���N�:*��hP6R��c�\G����uzX�g	��U��+Q��>~�ѡ$��=��/A�hJ�K�Ws�H�S����$�D,��vjs����o�huۥ/}�S�n�!r�QP\ϳ��)[ŋ�'8O���+-ܖ��%�*�E�<M}t���N�Xz�O4��	X2���Un��iҨ}�x��xNF� I���[�<�i�%��p/��Z#���rJ`O}P>i�͎��4��p���[
ގ�J�?�*��Q����m�GG�dkO7�d�|#j���ic�"��o!4.}5C5����޼���R�"_ e�RI_V$7��K��-!ͦP�����*�����
��:ᣲ2q��M!`ʟa7T�	}7���Ej�.8.�(��~FN��Dq�hYA��̋a:)<!�6��ZZ"13z3��7+��h�4bXI�E���8F�" 0�1���� �^jn�4�u!S ^<,U�H��υ5�������Q�>VNi�G0�b��6yE8%j����,��k8���2�I�flƋ�_�i��Y��R�|�A�řT�_*Az`��u�2fP�	$t]�!\�q	dV+@�`�BUV��<����?X��#�\��sd�ٜ�AI�9��a�͌��im?�6��x�a�`�,NJJO����maC���P���} W�JԈRwB���)��BbL�m�7��=�A��q}�/�f<�v�$��ۄ���g��#z��a����o��|�4�+5��	��X�ݔ�	���3_?	���܉�kRa�ps�X�����z4�j�u�^��J$��c	�ʽ���A�Y��tV�+�|R� h@*A(�^� �գ�Ǹob�v�WRx:r�R���G�@���]���>m 7?I7̕��[*�:�D���ˮ۔��6M?�+�~��(��>XB5�{��ol�oQk���>�yLzwxi�Z�ٞ��yCsG�'k5I{��4�O�#U��bН�Cr	p�t_�T�s�«�6�܇�_�¶|��-|j�Ln��|���1f��:�X(�)��+Y̋ Qa:7ϯ]�+o�8��>_��J1w�A� �S�u��tj�nQ@����o����t#��H�+�3�̪`��m�אc��R����a��)Oe>?U�f���b�2�{9����ɕCC����b+�l�:���c[�b�߁4"0U�Д:Z�mg��p�;������_�&a�Qvuۨx(�� }���V��Y�G�������wh�`���K�躵�
̠��a!$�:-��E��}��x�5G���t�
�^h�z�HO��`�\~���)ߔ�IS&�*��񬩥=_�o�K�T3��Y`�O������7ē�䆈BN�Q�>��`�9
�5�Ҧ���T2���bgN4b�'�,�W
#�L]����喙��c�&v�Z{�]�k�Y��;9Mц>�;�\<�MR�U��g�E��H��D��A��JF�SU#�T����:amuE���q��j��m?�##�^	DþJXz,�@��-�Lam�F�zR��HB�x���j���J�!��As��z�l�~����BW'@Ԛ�v�B�~�b��v��8�E$�nز�7�x��ͥȢ�/.V;�C�����^�{��߿\ݭRH�,�q-�\s[���#�<]79�U)�=m�u�A�>#�®4m�A��Ƌ����&J5�Y�ܛ���h}�t^e1�����k�������O���@)�T�cr�baΥ[�n����#�����Q�KwNr�9�FȂS�
���]����8ɍ��&�h%�
^���*Ff�I���Zf~��t�dqՂ��x�r�-O�~ HI`73R+�;vQ���Y���7��f�aBY��
l&pV�~6@=g����h��RB��f�v.)�-��6�HR/�ld�$��Aй�l�닠;<D�FǤ֖w�>+����*�+9#��zR�i0$�H���_
����T����Jg��`��d��Ȩf�up�&��=��h��e~�D��q�\.��LA�jU�k���#(ka�vR �tf�)(����=�Y,fq/��XC�w�np&����j�,&X.��Q�fۇ*�rm?�n�k��l�qOk	9e�^�HvF hR�����Su2&��*��gu�G��+���V�	�g'.���� ��M�YM�,d�A؁P���{�&���@aV���4�|eh���k��մ,�Jw`�5��oW�#2MnY`��ϦE[���#�g��(Z��j�X�+р�<�b6����ϯ�p�0�B?A<�E���ؕPY3�4��l V��J�s�檡����(�{#��sQ9����V@dsZl��9eZ鵌R��Y�\u��Ȋ�/T�����yHե��_��}���WT�-T-�J��i�wy�8��6��u]�Μ?������Z4������´��Sw�/+$lЙ1�{�t˿�RF)?]tnW]9����ޝ��>j"��F(Z��ߐ�9��Mô��ʚ�my$�V	J_.DK��d�6�sUMDLrl�1{�Cэ��
Լ��[RE��-A6�ȵ�DGA%?ITCW�� �^�(�σ���E�����n]�ŕj��$���c�y������f�:���6�W���9v�7b�7S�y����6�L��Z>l��)��Yl�]������3�%w~��N�oHR*��������cK�SyiT��_�����i�ɕ�3��	ݬmI�:���i���$K��束�<��źM�.-|��ΐl����ۀ6+�;�i�]1�FO\����	�&����ś�-��%�	0�^7��<�|��Y�t:�ݥtr����8?���hMvKy�ǓV9��y6��S�����F(|G��#���AI���N����!JQ0�<�D�G8f�b㛂�c<T�p�.6�O�#|V�E>�s{�u�!��F��M�=�+dR�$�}��oح�Pe��eV\�s��|��%8��@��x�c�D�ѝ�q_Lt��|� �Ul�15En�c�JHS&$�c�=�^]��95���Y�����b��P���$�L'U4k.f�ǣ@2H��3��������`��aK�j>��ό�{��hK��?�ٱ���2TL�̼��-�z�?�q
l^�#�l[q:.R�V�5�����ρ@�~�����.�eh  y�80��!|Yh�
����Ƀc����Ea�]H��$6�TzSQ�P7��;c���=����=}}}j�Ѩd�ƛ-��*IQ_�t6�.����M�-\���2��
[���J8��٬����֮���*^�n��w���ໆ'�n��lo�°o��e���FŶ��Qh���o�����K��U4��d���w�7D����;-9�uւ�;*��Z�3G�H���:���P���,���^`��' ���
ަ�	��P��XH㬢�=p�(3̘����asuX*���6s���{8�!�E[�X����y:7�X���Ub {h�Jm���B��`ҍv�ˣ\�*�C�6�_n�%��[�@�{Y�H�|����c�y�@��J��!Jvj�I(���k����vC���ط�X��LXg��	�F�dL��䝏�CH��l�dX�J�ބL6JuE�R�ߏ8�{78}�1��Q����}KRGS
��.��F�m��*�����͚x�-�
XKA"�=y���a'���q�����rhBaq��-��;��[�:2�L���c�f+iGxp�ðc$ܰ��:��^I�O)�2�@�7(�]�G"��`�6֮V3<p�Dm[�S��$�̨&���͍?�h �`�������9�|�P����M]A߫�g��`���3ʴ],7[Y%�s.����%�ؔ��7Q��������$�m���돋���X�GH�p1��9�^����?_��X΀޲M���B���
�E���u�����QO/:�����ߔ�F8שo�dLPc�L�O�`�r{���w�nZ�{�O��A�� �X���`�TZ����ۚ���)�`d�A���Mc�c���Mc��߃�0UdO4<��3[�C��2�h�vRY:��H}m���a��iO.V7`��D��,�ZenIL��Ȟ�"��H/%��:0�����,8?��r���؇f�}P��Ю����H�����Z/\c�� #������vfJ�c�����N���L���إᗘ�v+˞�+�J<�C�1%񪧓Y�V��B^�ҟ�SI�i�]�GM+,!�U;�8�*Rm�
���:L"�4�����*r��hu���t���`-1z�E��-:d�����8��ʓ@d�d9��l� x�y��2GGH�	�1Xj�
G���'�GE� ��H}(����*8�2�^�+�����Nه2��ڲ�s�e���-�+��@��P-0��X^�� }�i�0[��1�MB��שׂ�%���%B�ѡv�J<~M`S��j��<ύ1Ύ�t�����iv3K(z�= n��r�i���O������g�4���I��s^�
=N��E,(5S�p:���P�޷i�!~�z5l2�_>-�BZ�q��(���%AX������Ol����#fB�z�^�x담O�<��D�|�.J���z:.]J�o���>��_� �'��Zz��Av~�# �8�¡�˲��R#��u:��q�2�_R���A�e�u�k�����y�~h�7�ZO�f�I��b	`h0a0�H�֤Q�zK��-�=�P����vK�]���&�3����ǜ�L�D���\y���t��Q�"5��ߙ���V�$�O�H��/~'#�S6��|�}P�чJӝ�L(�[�;{��⊇<�(��f#*����02w��yY��ũ�}h�Q��y�<7i�"��6�X�㫬����US:��Hx)���Q;;�Ŋ��az@�2J�֧��pދ|x��4f^V8�G�p�K}���~�j�DQD���<%վ�~0�*����ox�H�V)"�����������ڹL��s+�Z�ve�أO���Q:�m9E#��`�O�؏��r�|�D�%��(���(���w�9D�'m̩Dh��'� �������ܥ�ٴ��v������g�d�2nB���xV���$
�D��NS_�55��W!�Eы#�T��e1���f�4p�ʎ�oyf���N8�!���^� 
k��(�D/n\�{�Gb�"�'u��l���<"�<L�A	�ϗ���h�ԕ��I�+N�-��a�������',isX�-RmQ;�9H�y>��bWm+	ّ9�����"4�5 ـ��=1?v��p�+`p}J!���V�����ۢ;%'��Y����ohޓ�N��o7��|r =���"|,�����_�I���d�0�����O{S�r
��t9��-�ktp1�e	��+u< K
�@���⸢ח�.�W#U�.����M��x[jP[�����P)�� ~�P�G�1�eAe��B������<s�	֘�+�6�LT5L�2eA��Φ#�L��x.qeH�VJ�d�@�H���%H��`��j^'2�6��g�/=;��$��E}��S����PR
�n7a�@Ya**�@;o	��mzp��΢�{J��f��_t3��V(��2e��<[�@��m6��Q�ݴ��&H!Ni�����ZF����O���$q��,dR3�{ho3�G�9��\,v�AA�v���Xh>�NI�\T������ե]L�3��~��<�clV�����Hd�P��Y��<�����{ﴱ����k|[�t��=�A%�)h�s���p�y���V�Aڲw�蝌��P�������).�ֶݧ�xjM�B,�NL?�>|��hM�����j���F��ٹ��E�	/��W��(���pvK��=�^e���h�5�ʍH��hOf��x��beע|��	��]Rv���z��e����oG�����)�+�� _n-�wW�}�*�9l�ۙ��>C��@�6�|�~��! �c����� �uy]v��=�7@�N$W���ؙ���О~x5H��ʫ�T���|�ؤ7����-���m�gX	8V�'��pT�*w��Q�n�u� �AD@�Yp/�v����.w�Wi���KI3�[�Y��Q�/Fe
R��*_���)Zo�2�����G;ax=	.C���1
j�2��H��*�*��^�2�,b̳X
4wb����&��#6uMNQ�����Mz�U��wX��q����9����>-��u�j�UaW2)p�zd��/�N���f\�t�d���s���s���� IC|D0��|a�⃑�9���tmg���Oھ��Lͻ�z꼑C���_A�΁��*�8Y���U	+Lto<�e�_�Y����ڔ���3E*Ր?��!�^r9Ǹ8lWe�E�'B��}�@;�2�&���Y@$�u~ e^����d�W;��x���i�I~No��5���;�6:�bm+��!`�����,!��'A�q���J�P�}�mV���T�sս�ͱ����u� �k��'7�F�jk�4�z��T�wZor��z��#z�)��'3k9;�^��^�P�;�������4�d�p�I��U/� ��Rù1b�O��^��d,�9�����Ci�^�E`��z�)��,UB�j̭�>�g[�\,�׽f�|9��pJW��x���\q��\C�K���w����W+c2�T�Օb��z8�7��g���/�#6���U�P��}��D�˗!��r����80ȧ^� ����GG�6��%&�Ղ�� ��=d�X�r\���6UN.&�!��7�BU��<�2`�Ѧ0`u��^�]�Ȭ�ps{�b~��k)���$y��'��A��GʧphIC�`�1Rﾒ���yv���#���9Q�5�ږ{��������S	T�o�-׋��{'0��[RF�l����E�G��s�Ɉ��7���*�;A� �3��T����
0�ɧ��ޢ�$��!Z�ʥ�_�@�K�*c�zݡ���%U!fx��A)��ŉ��j�5���o,'W��mBh�F�Ìh�s�@��1��M���K�F��W�������:�����J��2��K`�_�'9�vM�Y�e`��&vR����ShE�9��J�<em8q}�ݞ:����~l���>������>;C	8��v��)�_z�����z�Q�+�.2Z����XG�m:�L�2����b�������F�e��.Ai��@3L��z�w`=PB�8e/�۰(�P���������#�#�(��c�k�%���,�{�{�5�Kh����S�滼��8�
t�gcQ�@�����my�?��/��J	��V��٢�g�#[.�V�20᩠ ׇ�Ұ��]����Y|-%�5_싉baݞM"&?`I�m�Y#��Y���nL��T��_:'�Y�9CB��|p�]�UI�[�I{}�K-\��=��O�%�وpf�F�V`�G|j�Ҍ#I,��IMX���]ȫ�/W��6�2�g��	
N:zx��i{�[����#����ы��)6(QVE<X�ی��N������r>�ל5ƕ%��� ZܻE��£t�#�["���ۦն|/�#��F�M�����]��	j�C��/M/�����kj�yN�Ca)��u�u���;��b�x�%�*RQr�_G(�4���c������Hs�A�q��6T)����/*�%,u�Y]&N�eW�DW�Y�p�%y�N�r,L��*J�*���D(c�<	D!�DA����\�Q0v��8O"K�O|��0y��z�Ev�Z��0
aں�V���'������7WU�r`�3S�Y(�x��/@���~�V���>���%������gq��+��0\��M55.��>p���N8�r|�l<Xs
RN�!��8ۧ|���Y���ʸ�@};���Y�0�x�b��"a�9q'(�A;%닔�զ~���7�~j��ϫ�YJxE���l��/��=h��vy���ټ)F�/)���x���'4�U�%*x����M��5^P��s?f��l���@��Z���17Wc�������9�jO@cL�"2R3%7-KgRi[���z��m�~a�F�o[F��]��iZ+Rj����u�s$�1�T��+^�Nb��sŵ��o�vh�z�~p������O��>r�#�\+'�5�w���@�،��ՙ�Kb�	p�(���8���Q�X�R�f$�"��ǣW_�G�6�l��֛�Ҹ�%��	�9���<��:��aq�/j
u�{�c��B�_.jO�|o��j��R�L���;���3Ƕ�<?ђ��2ޜ���VQ�C;�!��oV���)0���ϰ��5r�A�և`5� ��ڇk�_H�c�%#����;t�	ͬa�@�	,�Hq=o;}��N���Z0��a��X]�QW�s��}�-�V�"�l����{��Y�/;��q~�@(w��L�Aӱ��X�U "z����B�-'�����(���+����(�S�_�vZnD��5sw}��ݬ��|?5d�����oa{v�|��ڽ��ԢE���CՃ�Y��޹TJ�S~�Qk�O ~[�����r���u�uSNLrļ`���|�����J�7����I���5E�P_t|�u�|_�#��	(��0�P~��x(��p�;�31j���Y�x�7eN����u�#����_G����a��S����������aq4�T$|S'�\Ot�Z�����.�,�g<�����b�Q����W�l^צ&�__M�i+zn�X��t�X�Tc�D�����!rI�[z��q��br�<l.��$I�s�"�O��z��xK?�h|�A	K&
ћ3Q���]�Q�c��{�q[Z?�3�NT(�MFhl� �9�<IN����%*��R��e�S�f�VSO����9՜�v�H�%fz��Y�>�k4��ʲ�9o�\1�86t�-4�E:��3]h���B	إ�2��J�s+�/�� ���ڧFC��=�=X�\|�u�p9�t��N}��ΐ���T�C�.��IZ`Y}�>g&�����ԧ�"������L�IsA���x��Hg��C(<�Jq����.n݂iq>UZ��0�I=��KO(��>��0��9�Q-ٟT�D�ӛDa*�77gt1)�іX���$�t��c������s���6`�>���d&"z|��h��;�p��5P})q�2|�2��Ȭ�4�yP�;��*���r���4�<�V� ��9�a�� �ƴvjs��Ǽ��5]X6�"�x��'��b_���D�x�V�П�>�;qf=W3�k)�A�SPX~|glXQ	��$�P�ż��{�jk��?��ϡ�L��/Ұry��5¾�q]��3�w�|(Z�0"|�v�|�V�FZ�|������3�5��:�Qm�8���~b݃׃�
C/��SOؐ5>cܩ�T0�t��p��z�/��ֆY����d�9X0���6w6�,��1�������}`| ��T���=k��G�2]y�0�м��.��O�<���"�4��t�L��������D�$��dF�1���r�jK�L��bl�N��f���m�[#f��>E�D��\�~6ĭ�9񷚸��Z��C��m��|_�������~����Y�8-��H���E��8���:
��o��D_؏��ܚ���]��r��m����8���w�7��.�Y�VN�Z�,��]�>���7�b�I�_�;�:Ll�/�u �J?��)s��0l�R{6}�ꯤP�`�|e�'9A�5�E/f�5
J���"*w�Pq�ǹ�!) "�J�-�U�prID*Y����͑�
C}�8^mwŚ�s��|Yє�<�_�.)&a@E�V��Һ���N���փ�ac>A�s�Nr�8e����yRH��`���F��=t �$��;e~/��V�$ZW���$��
ٙ��.���$0�Ȋ���87TV?N͚��>�r#Ќ�~+Q��Dy,�k���捖��D�Ϲ��s!��f����F��4��8�$*�w�rE�Q�O�o"����\��2���]$=;
����4�v,���I�A{�+���`�{�`v+xP�h�s��1&}y��'!��w��3{��2[������?)y~�.�=A��t70�'K��6e�%���B�H@��OB]l��8W����ؕ����O`�gJ!o?�%�LV*�i�^��!�͝��;q���Bj�������J�2p�O�.,����pNJ0��A4��
���BP3uցO5p)���˚�I�^����f�xTN�Mq<M21�ʦ�r��R��7�r\*�{��/�F�[� 5�xyB�l���۬��f�9�NI��V���{�s��%��ھa�[;1����D���M�հ�,�\�ŊV}�:A�c�a�,0 �7hH���f��ۄ�,c�H�/���u����9H�6�X�7� t	�q�VM:�T\���9kb��+	?P?��K��b���4T'�����'W�}ٮ�鸑����{�dk͂4��쁹�t���2�-�p��O�L�������a.sp=�_��ˢ�
(7�}�����W��0��X@)�i��ϟ� 6
K�_{���K�N�0��0t��A���'�q�m5�b"�X�jڣZ����7�u��3��v�֍�F/]�ە>��W�$����P����&/L�a��
os�5�@B�4}�r8���]3K�P��G*�$2���T��v���z�O��-FL��aN�{R��$�o#�p͎��sFI]���Mg�ѯ�f���X`�1��.ʭu�0r��aXF8��	�H|�l����@@3�3zy�D�^Q���Cgr�6`{�
���S�T`�ʞ��L����.��mD�7R%M��/fW&��ǳ���P(�{4�o�G�۞�0 ���|"�2�G����9�C^[�,�6�1��(�Z~׆W�#-s"~0������I���6P�оa�|6�-'>��L�����F��I'ǐ�*-�,uaa�uOZ������_����I�n��U��/��33��Y�J�t�P%{�L}��0H(��R��d�⣇��=ZXT�}���_�UJϼ���8�`$�^�7-�א�����$S%��t^���C�]�¼1�b��k�,��\^Ѡ�5I=:3�F'L�"t:_B�e6�w{H����K����?��4��J]z�K�X5��w��.8:��%(�eN��Ȑ��k9x��;�dA�U�DX*�2&7F�:,� �^'vQ�%+	�&�eO�;,Hs6G
�҂��s���1���o4PZ��*Q��R7�mM�aō{��W���&������Ktr����D�y�C@���-�H���w5���zr��Ae�o�f�jUE���[$�I；����U��Kf�`���H�b�- 7\.�6#�9�<S�
W��� ��2o�w�ɍam1?DX\��"�v�b<:1r i*!"�q�8���4���,�$:�4^Xn�0� $:���w���A��`hPõ�:��J�pt���͛ڳ#�tZ���X�K΢O��i$y�d�@|���ȭW����`�f��V�S~���v�xzX�˺�w�������f���/�gCm��3ˤxLnP�d�
s�2�{�_���0����q������'J>�;�`�0��
�_��d �v�W'�@`��]�H!��TR����[�#���Xj{���Y�BH�|���a�V���J킀�qݶ�<�6��@���:w��_�e���Ƞ��!7�,��+�Boj}U{��F:`�'��������j�Pv�k<��3c�(�TB֐,ߍR�d@�{$����i�ڵ;���6]�������yI��kkJC�x^�:^��	>��-��iJL5z�U>"�ҶG@�/�-O0V��+^ ���S�c�Ru@xI��;�_CkH����˼�l)�y>%,1��2��Cvh6�'�e)G$�4����B/������d�����ٕ����7a�W}ѥ����IK�D��O�a��_ �.4a��Z ,{԰�L:}���*i-?�p�G��k�P�#�X���	d�t}�刱oi��ħ�P�a�)	:%U��ܮ��/$,�ɜ��X�B�y��g�\����)�&�Vl^]���$�٪�����F���WG�*�5]�(���wtaw�h�S���S�6���ʾ���/f��;�`���ѧ��y��
1���uN���ݞ�b>���G.S�6Ԑt�[.)bg�u�j�Y���V*T��F-T"���-��V�6�L�g�>����^V��I$P��Fsr���L7�0��1��~bP���=8m��qҤ
�B�+'�+t�ȼ�wp&�*��}�T��Ӣ�,��\sVn�e�_UU0�W�j�1�̼�ӻvZ�_�g���&�*\�޿N�f���ɱ�����
Jc_m�D��܌�ں��b��'P>w ���jK��/���)���u,����&����U�r��WW��7T��.�������zw��Q�(E�ֱY����c��E��z�Upu� �VؿmY9 ȵ��m��+QV"�6�ru}8��O��ۖi'��I�>�V�cLh}腬<�;%�^YØԛ�zW>��
y�S�}5Mi�w��V���n�H4=*��L�*4ԇ}B@D�#pS���_/�Gf�4�:�@��qD��o#kXu.������p�AFdq� n��e9%������E*�Y-+���1:�Y]
>�xu@(��-�"��}�yL���}W�x�V��>뉂f���N�P�b��l�V��-�"�� ��e�5�M�ޤ�E<*���P��P���-3�9�o�<�>�˲�����⻀5"G�^�����7*��R����v�,���M�|6�0^iB����Ħ�c�k�p�Y���4V>ʍH3D���+�Qz�'���
gZ��]�gd�ȧ�����	#������#g�}+຤�
Ȁ�`*���̍FՅ��LМQ� ���Y���Qs�jx�J��?��\Pf0��	c,���F���r����ց��ť��{�ͷ����?���RF�u��|�dZA��u-�n{|BD���#׆ʊ��K�&����r�\b��Am��D�i����I�KڛWa��xW�D�w�D�m^&�C/e2j4V��	W�Ƌs=��K,�5.)sa�4@>������l����Qf�dHo6����id&��I���E�QҝH�T�[@!H�,��{���Y�v��O��~a��C�m�y�`��V!&�o�Šy".\V9Ř�)��_^^{3����	|N��\�l�o5'���NI�uɵ^���FVfȂ���5�>�� 5!�A�9Cy�~/�����	�E�@��Sb@���\*]A���[�M�%ݬjt����>�<�Q���cpfg��9cہ�dW H�8�G��41��Po��%7jȩ��M��I�՜=w���8��-+8��W�4��� ��E$P�>��*h�A���������W,b��/��D�Mc���
4�S�#T2mlc�i.�q�v�To�B��W��i��r�dD���tR�β�a�A�,�g�3۫L��ԲD�Jnӵ��O[�ʛE��E߶/�E�������l�T�����\|����0 ��2a���'�ث�D��cdߋ�ן�Y�V�˿M~�<�Ռ"���� {2$j�39%k���	���U�� �	�|�B��(�w1�Mr���K�'�*��C�:Ռ&��o��@�@��:����2���'9��EQ!�%�n�07�rBF���r׿� �K;ˑz����WyV�Ο��F��(i�V�%j��l�:J�;/�O"����)�YHk̝���ke���L�A��Q/`��nTRs��֭�����ӳ8��������ZQ+��
��f���\��j
'p�V-W6���HiI�R���z(堟 ��p�[%��D�*w�}��ӓ-�F~�&������D5�[�LiN�h��^�����w+���=w�e�M}��!o�#/jPǣ���|"�*=�/��e�)��ɡ"�f�*�s�Ի}�űΣ����e��Bϟet�a6�mք�y�O��g��:'ˋB�0��M`�l� �S��Ժh?���be�ר�*k�6W��qC�pR- �3��?�<�l�{[H^f�6`�>�R�DgxBJ��K�Uɦ�i�D��I��㴤_���a��s�.�\A4	��*zk+P���D�C�h�J�s��dA�㍞����\j�|�M~P��h/�塚x�f5{~�T�U�����͉��7�Jֱ�@����d�o�5:��v��	w����K�5O�>y�
�v�ҕ|1%��X��1�Ճn[���Q�l"!l�A)�O�D~�(*C<�9�q�K)�a���,�LɛNH���\:���$Ae��c�=c�l�֤����+�Хm�|8�J)'K�`
^��&��'���EE?��Ł=��]}��$~u��(��>�D���x�G����`l�@ŷz׮�D�v���l��v�ۉ�/y ��tk!0r`	U8���o��C��J�V���L�1���� ��U�g
(ڼ=&C$nr`�O�*>�j!C�ͳ�0����E�]V�M���ᬸn]�8�7�tė�U�����w�, Z�܉~uq��O�})���D%���!7a(�pc�q�9��8ފ�vE	Y͵{���Fx��&�>]FdjV��h�7j#`Q,C�B| �;��I w�W�uI5Z?�;e�7o��r���)�e4["�W�<髆s�D�踀o�dGܳ����z��2U�z���X���'���HC��5�"�]��S/�Sm������[���n^h���Gb&���{r=���޽�8"u���Z��h(���C�~͐e^�zũ9�r����������ܷN�ϧ���_!�	@$�x���~J?�'j�-	�TH�z���������i���t��TþC�ᘱ�3��p_u;�'��Bf�m����7��Dv0��l���ޔǧ���p�S��0-�<���Bg���:�dd�y	k,�e�[튍W�Lp��+�&|A(�
m�JG�ynL�Ү�2�@�Of�&��S8�E��2�4Q��p�6 / ��"p(��]/R�^��:2o����:�_�C�,=m@�s�7��̢"m��!3-+�8��jxh˛a�Z� ����������V��>�`&�[=w��C%���ŗ��\�e��i�ڈh$.t�I`���Q����!�����>��d��v�s.4�%���|��B2B�(˅dĕ.�q�m1�?�^i��v����_oyj�*wZS'˽������h/���~�R#Ń��+=[8�7�kĂ��y��T��>����g���Q�s6�֫�]܆z��f @,��~��Y�訢]�h�UWšxPp&V,r\Bj���!�T���4ߵ��T�Θ��E�s�����������So�f%ɖOc-��m&��O�`6�o�6H����A.q����p�d��O�ΝVO�Uy�
6�,H����!��~���_{$�O�cԿ���_�I�>�\�K��s��i�y���H cjcS�>o��Ə�&WҞ��Z��6�c�MA�w��J�E�٩�V6cQ[G�&�H>h����w+g_�8���4j�r>�x�T��pX �ލ�jɁ4�V�����`+�"���ՋL�� ������i�`?���K����AK3j�\~PM�k[Ù;��B���?�@9�$dJJ&TP��+�Ӧ��Y��S��]������N�	}��[y���TD�S/^t�h[2�iBv��n
����t�R�f�dX����X��㉯g�b�cK�g��ϼ���i�P�S��Y��^��'96g���2���}$�6�^�i���8�iN��e��ض��5n,?�I��_�3�p��	O�<@���([^��x1��ey�m���CF���^���l��v-\`ۄ�4�����츸 �	��i��xUc����M���"�^�_��ܒ���QH���F���ɘ+նA8�~����_�-ESFލr�;��pݨ��ޘ������?쨮�A_�}����jr:���r�RC1�$`e���='B@�̩d�{�w��jex�*<rY�i�/��.ǡ&$:U	0�k�f�x�^�}kĪ�'�1/��
2�#��`�5�M�1�	��bmw���{_�@K��.��z��\Ur<�7�d�~�Č�~����ɻ�| ����Z�`���@�4i4$	��U�U��\o�j�~��J�
��aE�C~9C�n��k�ÖBQ��	��!BK�Б��ұ�L�԰�ai��Ѧ��#Ki�����]2���j@��
k�@�՚Z��W4��Eq!�ء_�]��~��Tm��;����׵/5*�h��y����q�'�֞�|��0X'gd����c��(�Sr�8���V'4�+��g��P#��+$�P9G!D:$�r���}[Vr�*Nљ$�²G]x�j����I������Ҟ~m����񘂳C�bӅ���D���&���:��n� ��$�)���4���}�|i|��cu�3z,�1	��Oҹ�ON�N�� ��nK�< e&=�
�cT��	8ŭJD�
�H���A��wn���Kj���-��k�`]�����,O"��ɓ,d�rs�Pt���]����甂FErFt��X96$��9���� ��V�rEךB�Dϼ�/(���w�64?J ��"Z���s7ڱ�O:��0Xսj�(0ŽUp2{*��b�f�;)"�n�
LglK������|�@>��k� ��=?w�B�^p5O:Yu����M�"G ��ۚ[ �Н�-t����Z
k���<O�2=�l��<8�;� �4�`�� b&N�,[9����ҽ�-A�&����
��h�%\�M�E1���
��'�D��R�j6����:|T�ҍ�?�8�Ϗ�t@��iN�m2��B����"�+d�ͫ��;�w|�Nܮ!��Ga�u��Ovhuۆ����T���� l+Zش�4��[���}�Y���5�aaw��H7]{(�zz�he�G�2Q35�b��✻��ԁ��_�o:���ڎ�#�"Cj9��Wx.�{���Ǜ�����G/�>��&�
�{��#8�'0��L�k��]1��
��i�Q�͠�k�Z�k���t|������v+���ڟ����U�����T�9�si�ZQ�O��R$�o��	?i�4��� �<���������>�#�OM�����1�Ԉ�������G�9E��_�x�N-Yk*����Y3�c�m��ca��[�M ����D���N$~�A!�UUNK���A[�6W�������Ү�G�H9�q��z�E$����91�|��學ɬ��O�8T6*�v�4U:{27$(0Q��}S�����?c�O�~�i��wcK�(A^^߈�.��~6W _i�Wk��"���S�ܳiW�7�q�(��m7F��SnC� ���'��`�'7E�,3��URWO��X^�-��v�b��Ua��LTH	����j^ �F9�&����V��-<�8�(����� #��F�l��G	AU!�߻�,��aF��du�sx�� +^���f�L��{ê� ������;�}C�}�1M7�(��\�{�Y���V	=Olw��Ӏ��ԛL@��L7�	Dk�jcl"�h���CMI�C�7VR���^�^�e���3m+���u���gz�(�Vk��i(H��
��0�g��vdAp���$��#�u�#bqQ�'g���9�\-#�C6L鶍S�-�� ��@��"�sM3�.!nV|���>�
����V]�[��&����g�D�E���%���3E�a�]Y�h[�1`�a��I�=���� �8��g,#B`�y���e=����:<<��h�p-�
�Xc��>�v�����-�D���P�8Z��j|
���a���kP�A��O���Q\uE=l��	�������-I�4dǩ�#�ˮ��R�7����#w��&���Q}�f�k���@@�`�t�c��re]���<F][�7�W�md��.AwC#��t�T�n-���p�F!���'h��qr`��p~`}J}���������Ky�@����co?����U6eT�to� ���f��J������i����3D���z��)���[1���%�ȷF�����/B
@i\�Vq���=�N��R&�ڲ5�sU	�-I�ߥ/����u.*6�\'f����)��`��-D�=H�TG���ÉY1�n�_v0��w�(��R\�&깯���]ˎVJa�:�X����:*b����^t��4� .a�5�O��ˢ������~�·��Sh�e��W=�sf��u������2�u?�>�jJlCp΍�RC�@�D`��d�3�Ş��v�5��m,(G�C�և{ �|�hi��4��Ļ���m ԛ֚e��W�	a�5w�2'�Y��);�¼BV��e+ie�.�� M'�_ol�Vo�^�u�[�|���FrP�k4��~y>��ArPMW�71�v�p�D9u�H��srd^�����c�"0A�ܟ��\8�T�$��ۇ��Θ�Q���Y��+��#��:������Eش�rmf2�Om����-KN�]�X�!�!�J���0�b˕?�����)�ց�ЎZ�f{��g���#��=NS�����@�p+RD�x��o� _Y��mɹ�&8+;
��,4�7I���	ySOЙJ�" k/"�
1���_W�Qނ>��|�m�bu�xNOɋڄp���y��16,J
��b�* /X3�_铫 ��d�L��[X���:�
���V��DG��=��lF����|��a����X������fR���l^V��%7�S�y��ih>�@��⾰#�ni����ֻ�z���Ћe�
�G�0�e�����E��Î�7�?}d�;�?0k��O��\�k;����8�@D�-��?*�jz2^g���q�7���ʾ�����b���܄C܃��P�3xa�&���f�l��:��yi�(U�T%���F�O��ѧ�T"<�e�n
�����ƆHw~���b>�]<r�VR!,��qٵ"r���M�X��گY[17v���aE���5�\�0��6 Qq�L�c�ȓ�V���.�©�7�L�W�d����Z.�����6Ѭ�wT��(w�ׄk��iW���Om���v`
պ�A�����;��=Q��B����Q�h����q�?ޝ�|�u�]�x&��{QG���۫�npd��G	B��xrh����[�8%�������r��Ӂ��;���O�&�R��ڤ��i�������\ˇ�Y�<�qC�CL�܉@՜�x���$�?��[>��-KA�`�t���	�ɿHrF��D�@#���p�R ��tr�S�����x��x���T�.�A��e�@�h���q��fF#D�D1ѐ7������2��,�s��ĉ�Kn8�z$y��g$pKg�_[8�����_���1S}�N���dR�� ~�:X��;?)��Tu�� 8E���ٮ��~�魠�E^Nᇒ�y�7�@��'���#����r�wk�;�� ��i�FH��9�ǈE��bTm�3�6�Mo�l]�jhb�n6�a�@hO��in��+nrW�
=���s���9�|ϨK��]�<���X���A�R�Mmq}���~�Y��7�zQ�v��V��,�7�C)����b�zQ�w_b�q��B�ն�h�>�S��������6��9`��XhY|\�P��j�e?�}?�
��_�]g%��unx�����tęX��` ~c��ӕ	��ާX##]̣�!,��r�ۢ�}�H?�Fb�篱)@�xq�Lq�G�S0���X�<ڬhF�SyK{�Q���VH9AH=��&�>��O�a�ŝ
�MD�Z�K]Dk�c�w٪N����&1 	j?RU����F�K��ʷ8��A���n�ً�F�|z��vI�\�,',?Cu�=��/ϑ~{t�s*5Nݩf7-cgEQ_ugQi�-LG����40�Zn	���S ��Pޫ��~s��cf�w���X~�ozCO��߬������R����}�ak�\#:�|XB��l�d��b:�m�c���� QO*.#y�F~c�bO��e�U��+dVc��3���v��_�ُ{{b���bH��A������U����?�����z=s�Ȕ܆�J���<2�X�9���l�7��߅����%;���J3����St/�ԸA�[��@��"24?9�)x��6�����G��Uwԫ�r^�]����!0?yJe6��eMl�j���ﳹ���³�( ��U�/�����CA;VQ��(�2M�,A�D�3�#��7@�>�k/�ID>�w{a�Ő0$D�H��YsA˖�<�vW�؇>�@^z,'�s=�$2Q���{.�ƛ���牃����Ɯ���Tw�Z�Aqd�ɧ�@���C�u��7�f�?R��>s��z�����	�J�
��h��G��y9��VͶ!�*�=�fiǊ=~�j���`�҄%jV;����e!�M@�	�9�ۄf�MT�)��R���iC�h.�k?��x�5���=�֣����
	X�Ud�8,��$V<`��Sy�VL��F�����P���c���i��!99Q )(�1S����W�����4����(Uc	D��g��M�2(���1��� ��#
�8/�O��q|��p
h�n���2at-���kK����I�>�},��چ�nI\N�ea��Q4u�Tu��yl�f2Te~�y{@!Y�8hfe�@�I�G@ێ'�r{[¨�㤁�s]
�yȸ6QC����� g(�^�4w,*w���pb3� M��#��9�Q.x�(����2��S��+:�����h�)^y�HC�O���=��>��V����d��K��Aw�D6mO�8e���*@|�T� _V^����8�M�`�m�8��&
wM�M�1x�<]�)e��
۞8��a�	1�w�!�e� �q�f`XA?�4Q���⪵혻����/���z������F�y�Y佦yѷS��` ����Ù��|QǶ2�z���/J i��4/+�Ʀ����,��������w��x��Ile�15gn��������ځ�
��m���ɬ���%d(θsR�V'�>O���L��yX<?ѽs���0Vb�%TQA9((,(�j�NǼ��F��wG�+��<ZNK�ñ���7��%,
f��(R�el8*ca�y�k��<I��>����އ�ۡz*o�ÕYQ��#��<-)�C�>%l�B��հ�gO`F�+E��H\���;�ց�A��p��#_������˻����J�'�;A�[�>��j��;Qq���t��A���ie5ZSlW��n�S�C���.�;>t0��ŭ��lT~@����� _BVZ|)e��'ې���1c&,���!
�e@�f+�+���tD���F����"`D�����[/*lQg!�A���%9� ��2.X�w)��v�Ӕ��f�-<C�V�BP�ٗti��w�P��h����+e4K_���`J��8�QV�5���A� 3xkB�
�,W!��b������:�Y���7�]��֙�������������E-���Ҙ�Ʒb��%�q�r}⤦�yx�Bs���p���ݬ���p6\r��@Pϴ�u�$�ܭ�"�?8{�Z� ?����`��fB77���]@U���cʶ�V'�̿�n����3��B���MU�=�a�O��.3{��:epG�yu�,З�@+��[M<��c"6'��a
ˡ����A�VyH��wU��q@��j���,U�yb]�k->����X�A�2n��4R>�қ�V�e{sM���1?L�Y�c���zO	}��2��C%҉�A5z�+�V���o-��n��T��"]�E�z������i�0b�W������\&XА����(LR"1��D�vᮔp[d�hH�ʴ^�6�7��7��swJ4HhȁVLf
�]$7Y�'Y��,k(� ��n�p��m����J_�a��3��<a)�U>���7!o��O���������T�tC��^
�r�鿹�7s�?�ƥ�I>����Bu�*Q�O����P�V�(��E2w��^��f�m�H�$G��<�+=F�n��_��d 5���������\Ti�``X	i��������*�n�������]op�$A��8�<�nc��@�� �����b;�0��B��'>Z�@�	]֗_���`=���;g`���_��ܩ�ND�^x ��R���["&��V�0"��{Cht�!A�~�vh�n���������@��2��$}V�ӌ��9��)l��W��{���_�����#8��L��
z8�7�8.vR���1Ǜ�8Zк�Y-�;Z�|J�['�ڣk޻Jf�F 6@�Ĝ�u��v�	.z��p@z�:��K�9�\��R��[�W�.����;\Mp�Ӓ���
l]����2{H�/y���:V�
`W"t;��S�1-5���D���`p���w��W�`�fE��yN�#�F�F���c������x�[�����ǈ�X��yZ����YP}:%��A���H��y(s�+���*�Y��Ox�%�4o��� )�5�3\��ڐN�E����di&Mq���ml~P�Z�1�U�Ãf�R�}�P�?�]�����0ƥ���J�)�k�^2-m&h3�*i�o`��g�[�q_�����?k�[���a�`D���mney+«�=��и���E�����+uC�ڜ��-�B�*>Ĵ�ђ�}rv�ˍ���.�>[�8��hK�g�"���=��a�ө�~��.9��ʈ)2ǲV�i"Z2D�3CirE�ȴ,�e���@}��>g�����#�B�Ҫ���\��9�Ө���뛕AOO�h�n�[ԖZpe�=�z쪷�|��^*���.;��x�B�4�ժ�q]�G����[=`:�����@<Fv?��@~x��rYN6ż;�|V|�9�E�K�_�VM�ӽ�tS��7H���V�e
}�������}�W���y�*�\X�)D3�ޫя�qaV���PN���7X>�悄]�Q�:�5Saj�G�����@<��'�,�����ڰ��� k�S_��4��>l���_0ߝ$Ǵy�[j}ʬ,���#����NH�0f�ے+r�v�B��~{�[D�p�	��SØ��&3�p4�̳+���p��D��D׿R��VجR��N"��D'�8-xd��8U8G�B>v�`��P�����P�f������*�� �N����7�ʭt�)��$����9����FS7;��h�E�A-��&]�GN���W���v�ѿaG,����/yGs�G�����b��2�q$	�)�et�[�&��3��&�ty�A�]���r#� y���'*�R�6�PǪ�;s\?��E2�>��DQ+�^��5H����P�#���%!��^��%�b>vޥ�4V�CB?%�P��l�`|����6�4`�]]d�q�Zh�'�G��z^&�xf�!�h�<N�I�.4������# �I��y��tb��In�������I(�5���� Db�$_U����fvA�I(�35\��8[��f�&W�����ͽge^P���t��d�8��c���'��p��3}��7��������@� aѰsRY��-�ܴ���r�����Ǿ�7
���j��f�萝of�դƺ������?4�҅������+�\*:�LEf�a"-4H׽�A�j�I(���\�&��v]��mV���gۿ|�O��Ys ̻U��B����Q��#��ЭoK*���y��T���y`Y�?��T�ƍ�5�#d6�oS�耷�3���W�9�-���!�F�PE?�-�n�ُ�����`�Hel�=rNl�����j*ߣ������ �e�M�K�q�;����s��3�,*#g���ݼ��S���u^�A�M��Y�b�1nn{�o�/&��v�@0�nJ&v��<��^��N->v:���\=H*ӵ��a�;⯹u�*G7��I{����W��2?��a�;pSR>t��m.N\lp��q�js���o��8ڽ~1���b�K		�8� 
��k꩟��ͼ e�O���4E����|})]L�r��wFø��
v{�Fp>�,�O_!*�I�=J��J�I�F�}�tЁ����RMs�E�@�1^ ]+6k�Ǵ��d���v��vU�0ڳ�����<��dC�����9f��D�p�1�"�˫�^��`9
���p��#S^�n�,�ɦ�3܎�kj�.	Χ��U;�8��A��jC��DPo�Nʻ�!D� �[�W�^g}�03�J��lo�kez��H7,���T��8G�1P�@�U7�噡�
z).�u���WU�N|U����=��y9VU'���>;�ec�Q�=@*����#��q�wޝ��'���|]j����؆��7D�O4c���"D�����u.2[����~t�fc�Av*�rd�Iyy�~�����G�/����NJB-��bڃ�)4�j�T���੗z;�5#Z�V��H����d���	��p�Z��F(4�M��aG��k2b�LE|9LY$�������'1(���^�):��Q��\}{�P=����[��M�4�I)z{zLx6a&#RPy��b� Z��[eh�wY� �6
P�>�2���X*)檱���8����*aN�gu.YV�N�Pl��v�̑�b(~��<g�"]0sR�t;�,�`qy[*��8뫞ĮT֒>���a,�k�!z���3�8^�����MskV��8�|���@���Z�փ��6N�tƑJ�H2B�k��K�c���K��ip�,�
k3�9��%�ͻ���
��j��ؒ~'U>x�;��3>�W�_МPkjv���@p��K�qE��4�TP�ȠX��gvhmj���q�.�r�F���&d�uq�[��لף����8�W	��p �=WX㟤H�ƶ ~,���:3v?�K8��}����/�f�$�/�4���ϚmS����b���ҭ,
�5^�kv����|<P:ơ��z���7���~/�J�"O�����(�E���肠Z�`���5L��gS��~^#~��z洺S&�ޛ�_Hj�\l��t���0��w���⠷9�Ɵ�OS�U���aMK�yVN���e�OƆ"�:Z�{+o6���E��J�\���4OU��t�M��e���EZ6l�K )��E�Lf<9c��@+}3����{�[sA4�c�ms�þ���CA������g�O����Bb~,֯�S5�E��<u�b	+��hD0��� �O�?Q8�!zZ��}5��I�g;��U2�O���RR�G���{��Z�Z���gid5�=�IF�b�<q������\����.�z8���O�S�y|��&�v�iV�F2�#dU�*�<��x���cS�+ё��yf$���K;0VB#��F��"F����Y���(j�XĺdgAeOh�ң�]�}��&.�\E�vEarfW����~����Agw����^}2)6,h�v8�D�N\*�6y6gUA���i�{?8��f�̂f��xZ\���B�6�1c9�0���zoK���Z�obRe�Z_��gA���`1�� �����35�J��MQ��-1��p�NՓ[�-y����|6��ju�,	����~�.����8!n@�wK�Vq��>L��e;a
x`���0�(����O�~a�{�;�����UzkGQ���|fPb{�r��o�=��e����%����k08ѫ������X��p��o��q��/���+P����|�?k�N����g��� ����G���~Ab �4>Ew�^Aj�dt�w,*�T�q�Peї;��Ô��#�]6���:M5N�����1L ���ਆ��--�Rׯ�e�2w�Ӄm�.ǧ�ߌs��I *�R3:��V�]���P�&_r�xI0J�Ŗ>�e�_�@���P���C�F�����z��B�мR�.$�|��rF���w�:~�*d����q�V,&�����[��+���U���Էktr���!���b�z������@>�K	˥w�q����xIP�J*�u����^w��pԫ�X-���^�|�&���c�(G@᫹ݝE�j7]��ש	�ۜ��vӋ#�)��q������e[g04zx��A��R�l�@M0�!2>Z�092�n� h���T�����f�{��߲��Ct�����>�:;�#c��uȚ�Q�9}�KF�z���T��j��!�4�a��5�x	�h�R&�>���%��*P�M���DҎ��J��� ?����c�Nq��%�:{�����vj�񄘿��?�jV����Su=4!�Qǔ�1#�����-�I���SZ��$��~��bR/e���Gg�2�bb@F�*��d-Vy����6#n��:R���3��"z����k�ȕ�A�X�� V�$�B�i6�a�� u��M���{�M{ &�;�dӂ��A966�O{ ��9}��O5�et/ʥD�'S��MpҨ���Ld�5�ev��9��H�Wv��C�#V�Y���b������_�N=�� �gᨻr�uЂ��C�I�HT��lD�%'�����=z�u��G�O#�θ"F�+��3�p����\�C�빓��5�G��4/s|Vb�80���Q�����U��a΃�d�8@L���g����^�C݅y`��:�2�}H�A�� �<E~p*���9��n"�z��Jn��|$;�0�Q{~a��XhmV��%�@'�)�����fQvȡ/���������֗Iwm��.
V� JVb�q��؊0z-�ĪQ�ý&�:�Zb�r��Ҏ���G��p�}���
�_����>�;D��ɬi:3ܞ�'�(��y�Sq5�RO5n>��*Y��G�W�}�������fcᦄ-pW-]�%�w��}�~�N��V�`����|W*�v8s����yTh�Y2^8��lR�!-��T ��?*���f-��on�o�5�=)8�Π�YF(�>j��b�}�r�ͯ	���P��E�llk�>鏎'�&������n����}�?p����ɋ!�N�R�
@=���V{�]��{�0�����H+B3�\�O�K�Pn��(�G��������z��6�����p��da�m���Q���),
r*_�і{�ݏ�d`y��:A� q0J!�b7�.�T��:���1c4��rt���`�2��чR��}5M�%��u?��^�����T�DQqX@�� \n �q�8K8?�ʌۛ1�-���Ј���5�(�a4FN!�.�M�N�sP���d6�UU�\C�(�"9�jW0�w)E�V���w	�z�=�$Ȃ3�qQL�R�en�xV22Oo�K��-V�UaYo��- A�D�OGA��~/�jC�*�֤lD�U�r�o1Y@by�����c
����1�Wꛙ�	���x��<f.m���c�_�gB��صB�[Z0��b�+P�tͧ��}�?/Z���)�g}��3� x�kl��\z~ώ@ L�G`VU�v�'>l*"ښ�G���A��y�y�el���y�ڊ��4�ڎ�j"�f �T�̸p;���sT���}=�t���@��������M��ӵ+ԝ�E��d)#(.�OQ�TG"�hQ}��'	=B&��/6z��|��[:��D/�w���[%
a4	�+֤��S�ϸ< ��]�TtS�#YooQ���Q��.w$��1騥��4�D%��wu��Yx !#鶹Z�S��j�sV��pI�|��i��{��F"���k��H5/�\@�I�YK2�H:om�p���Ԫ�P��2��1܍LE���N-u�����C�ݠӥN�
Gɲ�f��k�$HSjD���*�G�6��ˡ�m��D{�9.�
*}f�I|�W�8���4@��Zֳ��U�^˘6;M#L�ŮCM�Ưݝw��a���A�9b!'��3�W�O���-c���ң�_P��-��h"��XΟ�xA{�G�m�	����Fq��{ ��7�]-�3
�K��欜����*�{�*�PV�N<)Yi3X=Ih����_A��)������u�l���M�z�_Gǋ#����U؃mCn�)��.Ib|��h�I酒�H��կef�o3h�8p���-w��d��/@g��,6��\�������0���9�@�X⶧��	\:؄zI͋g۬w�6H�7) �>��]�Z��.�}�)�4�&cV�H�`e��MY�7����z�3� �wpb�Y.���d��w4aJ�(�3G&Ԃ���h�?l����FY��SwP�Cby�<�&����d8�L�,3S������������{d`F�d׮T ���c�x�����R����Ҹ`�j�����/q���⾖5?m6��&�	��a�*-XI�3.~`�	�Cf��$�W�-+�,W������R������I�0�J��M�^s�sk�����k��Ty?l)�����"���$��4�v:�S�`��
���G��I�nw��Iٶ�s��-P�,���e�� �v��4$�Nb��s9J���:feH�EC���$���@��K!�hY=/r[Uް3�z+�4�'��l�mf�Lߥ�FS�3�)�����3�-T�!S��n7q5<�Yb�-\�� �21)�P�%�{4}�����s�NQ���"r�B����S!�2���s9�Xǣ�
Z��႓>DV!��|�� E(`�BI�z�隵hF���$�sRm�P�+Ks1���O�("��հ��=e<Ksӟ,~=�a r{>��y���i���Fym>����DrjLC�_��3 a}�T���ǌ�*�̲J� u�񜺷� �u��/8 �oV�V����f�<�[6���a�E)�Gc.&��	 �/��[��W)c9]oH�J��������UȌ�3[e��I��YkF��Y�g�89N8m��Ѻ�t�e+�uLSZ��{�9;�P��b,�[��L�1M�Q������O�4#Ll�af(P�(��e�l��X�RoM
zP
���Ofi�!B<��;��D�����9ݒ�%�-�*U�]�O7B�1�@[ܭ���2�4*6U�L��/��k�ځ�Ua1�&�ׅU���f�j���_���L��3�R+opj���\���l������@�̛��i���͕���t����<N�b����-��i9�ԔhI�:�>�hcq�e�;|������&d��J<����k�,DL�Y oU���cfߵ������rC^���5�n�b��.<� ��Y,��P�5d��Q�lge4M/ �
�]�E.�:��jP�8?H�U:.���	�Ŵ�ضL�0.A��Gv��Qc��b���E=9�|���A�2�;�U�i��o	���~�����-�Pt��t����L���,
,۶��J!���%�w�P�֩����}�Tw:P�
���4�cZX�O�ː���z3���̻],s�=��]�il4�k�\H+��z�U�|I@b���VY�qv��pX߇f�)x?��ا�����r��r�4}7��"Jd"o�"�o�B\L��@�NBbG��I�� �HN�o�ھ�|��="�p
D�H7ة�/�W����J��ώ�e ����
�Y��,{����\M�gVc`6!d�`%���k�R�>���>���T  [��c[!p)�߸��ĘS�a!F!�WCǛ�}�T�j�X�K,��8<���ot6&H�^HyD}�B���Q`J�0��5&N;;����-��o!J �{����n�!�"q�K�A϶K�矫z>�P��N�1��a�g�9��mP.^�dClc�p���};��gg{n�����"?�P���^�����xk��t�T�P��/A4-��4��>��Sl���1]Emiuw�9ʨ	Fg9���4��,3k`Ͼ����T��!7,��pd��X��8d���1y��*�t���ǻ0��.���v򩇅(����fJ�(�N~n^��-ۨ) �]�!�JT
�������eq)<.��#���
�� w��a3xI+A~����Ȋ񤓕J�����Yߣ��u���ΗU����[ ؒV�<6������鞖Z�5R�ʩ�� Rs�~��6:�+sp%Z�ùT��N22�\�y�7��;V�S���!��������$����q�=b�O?ټ�ב��RX�g@S�>��&��A6U�`d���/��V;0�gZE�\����,�%	��\�F�ܠ�V�A�)�ˑ�Q3�Hئf�2�s� �v�p�U.���<zkT-�_c�ε�AE���z���H�`�<QЍd��g"(4�uz"Ȁ��D��[��*�=XM�m`�]���j�}�XxUl����?ou�ܲ��y;(������-�W�J�P�i��aw�P9���*�/��n@l�S\��&{�N��u*�*5�joU$s�Me�s�=��������ߋN�\�X�Ø��[�s�3���E��<a�Ѳ�B��]��B��DL��Ƣ�������>5�A�>v�Չ��%ыC}��A9���I#S���Q��w*"FT�6h,Ber�����WZ����4T?!_�C)vԅ�$�&�.�b���SD��	g��.Ӭ|S���,{dD�Vo��)?} ���?�����<��}N#q�|��|����S3��bW�p��������i��3��P�2�-ϒ�H�=!�lF��G�IYe��o�Է��6���*먯�2UT���D<�
�� 8�kJ[�Y�5 ȷ?�2(<��;n��ô"���q�7�@DZ����<yγI�Cq��4PG�eO���ʩߍO�?�/?�\luv��-�gkS�$Af�b�؏����m�y\���5Uu8���_�Kս��-��c9��(
���R	�-��f�=#m<J3
�ݵ�ap�����t���2T?Xy؏J?7�@�Ҭ:D�/R�q ���?B����T���άU�j����L�h3CS�a��
��7�J�-���Re
�^ϖ�q� K,�{��3c�Pxj��JV�sB�R��P�;<�+��^��3����n$�L����|��J����� �/T���؈���j�=pΫ2BU�jY*�_�v�{[
�?�gX��f�Ki�ƒ�j��Ԟ�d>�HM=O'b��N���H��ӂ_�|�_�Zi�gH�8��y}C��>Rfx��
�F*9����>č����뜁�Mt�*?�nJX	�D��f�PM+�����|�p��_^9z4
C�HXǾ��ɖ�ZNJD����dC�� ����$��|F'X�硘�}YṫI~:U]I��pQ���rL6���c�3Es�fA�@���i?b'Z�^�ؖX4�4���|�v{����~G���U��6&���/��\�������*w�Ǝr��9�`�ͷ�TV���䡵Bv�3:�I��*��}���b,w0mp�[VGk�r��jm��1��*b�j�I����Nݬb�.�X��}py���F�V��$|²�Bb���[N�	�y��L^�����Gv�E���f������L�/"K�]�+l�f�4���کG9�D��;�Rނ��X��@���DT18�P��#,}�"�m�+O�:�d�3�p���:ձG5��7��\�>1'���`y��ݏ�;!�w>��|�,[��>�j�o<$~\��)��� };f�%�Aﯸ��&��]3���\7Y����Di�\��z!�V��.b'oA��5��� _u���'��X��8�!��hcGʺ��ܣRw]g��V:�=��h���_��_nN��B�KO!c����5��o8���I>����C&�N(��*o����ir9k	�Y�F��~v�_�"��T��, N#О�C2�\禮8�>&��� t�y����/���5��0ƺØۚ^n���x������I�^ڡ����I��$����h���0 ��� �����Y�'��
�1.ԐS�
�*�G�E��J��;~n�-�te�E�↚��1�Ve٣bV,-�sh6#\���]	���tɛ�pHV(�m�J��QƩ��i��A����D5��:��d,e!�"���S�W��8��'�Ҍih���A��+j��-'����{��9���,��ȩ��c^⋻���E��2�w�Y�����5rq#���t��b"h�/�*�rb���>*O���̰�xƿ�f�}�tW��]��Pe ^����[��9�;u;�%����iǋ���s���.�r�"��"U��4��`<�������������gc��?��́Pl�QW��2�Vp$�y�'��Z����1J�°8q
8�Zx����O�Ըf��`Mk
�ӛ�����u�CsH|I��d���I�Ã�ϴ|�Mfz�����r.���Q�)�/&�n�%���#���1�l��?"8a9^Ą�L�k����qlUE�^��d�#\�y��<{~�XF_������X�w�@�龒'�
��H���Q׽��9��:�'��KJ�2 ��.�`P*�2�F�R�7֐g�%��{��_��0@�p�o_ǃ^j Z�i�L��I��"�J�:�WM��~�0t_��;�$�'�ƻ�@
[�r�8s����'�������s���;��^�iF����A4�|@a;������玚�%��+���4Q�L�D k@��(�#�>`�c�	P��9S��� a@9��.���8Pjj���9^�X/�k}%���P�R��O%La���<���6�O&(� �<)�:���с"����VFԁ�o���1hJ,�Z�(
��>���HwN}��"ãw���"��1feH���iQ��'���8��9�ȿU��rWw�4�S�Jp�FW	_o�qj�tt��X5y���&�-@��M�Wd�Ľ�[p�U��7t2�!�3""م|�/�u��	��`������L�
��M�U} z6�J�H�>M�ʞ`U-�<1A���'DP���DGW����9��M�/~v�Ǝ��,� ��Nht�azc��D�0�?r<��0e��uH�L�×��A�X�>�����e��8��U�d����Z���i�$;bX�*���4W?��pD�0B��1D�*GR�a8&,]4�[=}�״�u��<����%���B�4��8���;;Kt�o5��W8�ա��kz��g oiA���^���!��s��ٲd=�c7�{������N6XeG�@�ۣ��M�Q�'�;j���u���]��d��h�G�n%'
�Ie%�n�zY]8�=Ε�)I��_j ����>�诺��#:mhu�K0�����A`_+�~���6ia���n�' ^қR��!`%�����epz_���ҒyF��?�1#G��|�!����'fb���0�.�_�b�����Թ{�Dp��^��ٵ�-蠩�p#��W�߫��K،�<�������%q��G��&M�ѳOR2�C�0���rx����a����j��2q�$��R���2�;�Ld4�ZθB�Qd1<B�(�pq���q�ݷ%�5r3��'���3����A��"$ۛ�ٛ��I���+Ǌu�VJv)��{Y�WV�(D�ԧQ�nBm������W_!6���<����	���Y�*v�����Ͱi&ѻ�X ��=Ip�p����z��&JeB�7�Y7�QY�c�s�um�`.�Sf���A�xlƃ�?�a����i�
e���>����uGX���~����cqH��6&����_GeIU�^x1�DW�E��\���M@��O�3�t:V�[�ڵ�ՓQ��M���J��A�my~2ϑ��ˌk��<56��p/{Pg-��{�{�hN���4�c������
J��q���+�nr�Y�����gQ"m��[ �\$�����������'����^�mZ&���#��<�iaW�~�K�}� pz���7t"u	CM���A�Vf ��"'���yS)�V�W�F|���21vTԃE*1�Ⱥ(mtD�ӏ�ip�i�@v:z]��b���vmm��� ��ψ�/5���	����B��@4]j�Y�f��0�d!8��1ƒ��ogt�g7�q=���@�)3YP��Ӫ�$������!/�2:�;�B��Z�$���M����-J�_0P=�Q�,��2�6q��r�l��P��63��jJbP�.,MT���Qz��LP 6~�9�DT�|z�Gg�j���b�$qL�ň`�w>��4�L��-�|μ�P��D�a~�3�,#��fa�g���~)�yO�qŎ� S�ū���U@��t�QV
��3d��s�������p�9T��:�&�#g�C��e���H B��_t�;x�G�̰���7W�u��{� � ��=�Wb��sm����&>VP�-K���>�~T�&J�F��TN�B�k��2�q�,aǔ3�!�V�������:ｬ�XӺ��O����;r7��f��n-+z����UjDL���$E����zH��є��$ؖ��zO��P\Yb)i�GaQ�r1Ԙ~~遽��
�)��١�����{[>ʶ��E�QV��5,Ž�C��b�%���-���� �y�O8��dA�׌���2
�h~Q���X�I�X\�Zo/E�����pA���2�#�{�ʲ����d+P:G��+%H������G��qG`���f��SG}�j�5^��YKp��V[�V�����`Q.��=X�֨�3�E�����PD�`�FW��%niƸ�m/��Z����g����$g瞜͇~dw+w�n�$D� W������m #�j�)�[���}&�k��.��T_����B�	�8j1��c*�]�
�P,�HGl��si��Q�j��賞\(�o�=b�bk��"�`d�j�ݱ�e���ؙ� �5��b^����4;ԅA�+=�����}'^��νAW*6b_��k6�C��Id���e��'��Y�$�H�.��^�q|���:,�Tc��!�?D\.~c2�&
�q���;�y0]���"���e%+�<e���_���S�"!���B3�1>(��kj�;U��3�@ %�EV��n��9"���$�����+�I�J0���x��k6��7b���`do�M�'3!U�q��I�^_��0`\T�l�M����� 	8MqIE�wW��+Z� -$� �KZ�q����8i ���-�����4��:�O�!���8#�(~���X��(��[�*�(�t����X�����:�b@,=2�X��h�6�v��-�����驪��?�pb��#&E�'���YΙ�����m�/�t��<C���� :T��L���5��Y�@�SbG����i�o����1�|�w]���J�Jұ\)�Mߨr�8B`d%LY�l�����<W�ꭊ��ݪ��\�Y�iɜ�J�;��r��ЊF ����>ȳO��>X2Q�l�������f���gsߘ��Q,ԡ��$)(z�eʮ�u��G�5--,��&p�p1Ѳ���M%�
ݝ	��	��B���1�!!�	��ei�Ic����J�IF�aj���P������v ��j!y�X"+�mV��S�
�2�g�C���ǚYŲ�@!-�I:����ICM-�'D�6댓�!R�d(���dy��F�$��fg���~��-�C2,T�, $zh&�	5�T� e�iy5=��0p?��	u0]�9��$Jj�O�ƋJ��|`��f��h[�/ph�օ9�~_�<����o�����J���������=�gP�-��' ��F-��+�o�s ��l�ĜD;!�4 ��-a!/�.�i�Jak����.Y�L�B#[�y>���{�	M������X�Gv9�;��$#�Ά��4�E���9\u�kŷWJN,z��b��C�ђ�y���=�4�����?�� LѼ:�k^a���Ν�d�16���\ �6�,n����$�/��}\���c��N�$1�c��#����ކhئ��KE:�&�v��$�ұ�$z�ep�Cv��@���!�$��zbʰР��dኚ8�_aj���ꯝ�9��#��i
v2�<��ƃy{zq�� ��=�_�7��F����׺���4h��B�@���T*�J儻��lq�����O�?�Z���M{{����b��ȭw���쁝�{}l�f�T���F ��bK�����[<���^�f���e��-MHz����h��iF�%V:}p	on̴�,S'o�e��7D��Q8����g#�C{֧9��6"&�2ΰ��IL��J��c�J���h��5£���e������_lC���f \��=�˫����ת����$G>��4_�78_�q�_3�`��c���䚜�=�d�^8���?@�_����mᦆ��͟�9���0ￎ�Zja��:3U[rc���B�T�@Jg^q��g�S�m�uo�J��M�k�xf��0�:�5�GW>đ-��&z�|�!�Fak=!x�s<��
R �_��������z�ߧN���tʙ��vx'7�໥0�:��[�� r������<@Y�P9�Y�i�*.-g��-�d�2�9�p\T�}������}Wr��l�f3��33d?�+Mr��2	~ �='�����Z=��r�H��A|�ɰ" A�E�ј٫x�%4�	�U�nߞ1=��\��K(�.aV���$_�(;��Mޡ��R�Ę.m�FZNeP8�ob�m�8���f����S�nM��G:����׽�1�",�{�j+�?b�!�n؏zV�RbUQ����)�����QE=����ȉͱ�	Fr=ӧz��v31���.P��h꽅]��P<��Ey����Eg�9���(���ar�#e(��,�XS��壁V��i��K����e4|��A
�EcH?q�?����;�sӗ�y��__
��Kq4ڗ�y[�Am{��m�@6F�E�b�6��7��4,���R���jX�Lx*\Mh.=&�Ƞ]�z�pJ��cpj��I~AΩ�'�4�����a!�a����Ԯ}՞��F�����?;�h-�*�@�gY��b��9$�g��B��u9�y�1p^8pU�� Y��=x�4��[�r91��Z��`��|�9��4��i/��<�џx'�����? �
�4p����< 8���IO�x��g�tX�\q�F�ǣw�tX`�q�LzcF��H�<ǹ|�r���z�}'�m�́N��އ��|Fx$`�(��"�n\?�>�O�Ăf��d�����(?GH��Q����� �ΏS��QR��.�Gx��I4'��HH��=�BC���9��z-y���l.����Ѭ�g�p�%~�p���8_�T�o�L�>��$�׆'���)1+�w�p�h�i��eQ��!��<���x���:�	=2	���y�;����sQ�� ��Be=y�$j��`�0=qx/Rm���V�=��2bi�)B_N��y�X^��k��z�!�,�qc������os��?����Ρ]�)�0�$&���܌�{�p|���:��U,�-.��H��5Q&'�a���-���*kt�y{��.�̺��aU�8�z�Ni ~Ml�5���i�F�B����O��&�`b��F��x�<@�/Me�<�1�*=�Xo��"I��>��k��2vo�����J�e���}������R��p�$φ�Of����52�(9�c{ѿ3u@�w��cA�4���,��O�Y�����K�g�|B7�����q���{DZ;��>���+_u�r0D����B#Џ��=��Q�5EO���D��]����Tw��q�����ӂ5�������<�g�j����M�J"�OI�=eI��3ѹ����S�G��d��QC�����؜�K�ɔ+=�$�D̡�IK��u?�%ѳ���k��q'sR��3��ܞ(Z �M&�-�k0�~���^9xZp���||s�9�\]�>��j-vRV��8�>�j�%�62�9�.XqI~'����d[���7���(��ճo(ӵ�, �n��\���l�g�L�z�z4�b`.��ۚ�Ӕ��n�<4���t�P�.�K��͗�C@�Q�*�@��o"&�x��\9�+�3$��"c�
H��.F��D�*u��ay�uCC����^���W�+?�� ������
04�d�\�P�����;�h���������+π�K�Vό�a��V�;�޷N�Z0@���
Gi�Ct��������	�z�Fh��!B��^/#4	0���dp�`Эp���iK|����^=:�Y �����\�H��u�9і|I�p���q����F����	zU.Ȉ�\U���A���cح�]�/ڙ$1�[�7}����}(eU6Ø:��0sd_�~�����g�_nc�������qJ��>��kİ)�\Rߚ�D"t���,"�����⾤� K�����d �#����$[0l�:p9� ־�+��c�k��p�:/�o�d�qUB�ũ{d?�E(�9�x8�Lv譍�s�-�!铞q����ا&�%����>���4޾>xq���_O>1Pj2?%�ZJ+�N��U��*6<_��mR��U�N!�(X�b�g��wk轖k��"��i���Z�%bx�n�dʻ�yW�F��$�ŕF������v�(Z)λn�1�|�9/�W��BZ��w�"�H���p�Ϥؠ�s�#���}���ƣ
��b�=kKT����תI>��:w���i�����N�t^�Y�G`5�|�Xx$��b��8�<�LXl����� h�����G��6�0��zU���:T�K3�P�nKv���l�I��5�9�Ƃg�U����{�|�C�$7��A��`d��%�Mn_�|��!�H�)����1]�/k�Ӿ�t�����4�RK^��9F{��l�����	�
2��S{��Zިr���b� SR1l�i������%Iۃ�嬈��t&N��a8tHӕk�x�!5S�����A����iJ�����	@E%���_Ş ��L�{.�5w�M��H�x��T���.m�m��P�7�4�K��K\+ݥ���J�8��7�|!�L�M�F����*���Q�+���������w�pVn�����$�0��0��W��,d�(�bԐ��HT��yKU��>@�(^l���ʭ|�'M�\L�c���/ǧ��o�Q�d���w�^�A� g�n�íה`�*���oEP1]I�;x�|��jK����/]e��8ԙ���׃�h��u�	,������������e���IkL{1V��~؎D�?.5�J�Q=΂�R�����R`��!���I=�z[���ó��d�8_@:c����\��D�P�v��V���dW��wdG���A$#)S�fG/�*G�,�nO>�[�&�V�E�eP�x���6������� �o������+����痣,�]����-*�~��P��z�͙@y�,!d�(��\��\]�3i1Z�hHMm��h��ꏻ%��OWgH�WViN�7Ծ�;�<��9w��j�5E�jқ:+uX#z��?G �y��du3�
�|A���"z��<��0�+L�����^�\:��"/5.@o��(Y7�vI?�k! �*<���f��C�E$'��,��_=G���;F/�m�/�Dj<�����Yz1����G2���Qj7�)���W��E3������XSnU�GW��d�~#H�=QY�ԡ��t��;�q��"c\UE��_�C7j�m����R-�h\:X2����g>%,�iM9�{݂Pk$�G�i��9�y�ߞ�6a��-!P��P*��]c��$xR��s#%n�L3ZӸ��u�$�O9e�>�� * 4ھ�c"������,}�챨A��M�� s	�#(q2)�1.��2:����fB5�p��d
͐��7��jz2�O{ξW
��NS�F��B��Eڨ�->y�Ƌ�I��E���Vk���9	8?!&����P�D���{m��Qi5|��@�i�Q����g�`��g�卷�IYN����ȁtiXhę�,W�1J%�J���!�p&�,�~˻�3)���
��`9z�ʕ��o�>6�1 l�Z�F.�#�ф�Zb����Z���O����P�?�4n���I�J飯���=;Z���?�C�h�D�v�z� ��/ I��l�G���0�������Y�������;��:�ǾY�+�S	�M�z~�67�`�����ή9�]�",���6�锉��|�=)f�Yru���}��4�B��O����T���O�7>�#׎��Ex��k]���/����p����PsP�A��VG+wuM��ڌ�2!E��>Vn�1ɬ���oD�Yf�S�-v�ooZu'�u�:RFi�G�4�$\N ���IU��+��.O5+I��^u��OQ��,WR��<��ѵ��Ĵ��t�0�K��(ˇ��>��J4��V�1�6��O{�Ro)��-l��wb��ok� |R0� ��-��g�]�$��+� �j%7䬃V�}�ڿ�a�C�Y�b5\'J����m�j�T%���,6��K���{���-Q�}�+W�\�bhNT�t�hZ:�v9P���(���ؒ������c�ʲ�4`�v(����ްF6ڼ�"�O��Z�*'��樂H �q��������cE�H�7lm`��N}޹�H�s��������x��ħ�^���n�lE(�����ҏM�{���s�sū�M�6F�"�7���?��u�M��җ�ɷU
��X���[��h�icʁ��p�m���[ ���"'e��8&#`AIQ��� �Hw<�y*@��w!��3�X�q	�D��
??���l�(���ww�3'Y��c���>��xb���L���S�0}K���s����:��8GM�1�}�����N1I�,}�V�߁���FP�5@�����䠺��(J<c4k�!����m]�t�1)W��;g�F�|����|��p�!��/L)4}I)�s�I"`dR�נ�O�\�2��Ϗ�y[S�jaX�G҆�rgΝ[�O���mB!x���ʢ_sNQ���u�{���7�Y���ʢ&N�,>/�ƨ^\>Ŧ�qy^�(F,�D�Z�m��ˑ�U��}f�[^�D(�����6�l�_=���q0\�^!�O��W��m�|�ʦ�ho��/ ��cpa3+*@d3�!�SH+�*"N�^ �N�<�����Jj���n�k���l�lrdƠr7�pR:)�"?4�q�s܁!P��3����%hX�F	�1� ���EP`N����#�����<��n.�4g�����׉�Ǔ��z~0�; �ŖS�LéfCm�v{�V{EJ]`������9���+��%hG�"�&��?� %��C��������RQ!UC�����k^��8"�ԧ�cd������
�����: �c�N����`�5[7�@���
�k�^����{��ӋS�>��[�	~�>�D�����ݞ�$�j2V��X&оl<�`A��\0�Pb�w��*K�߭���+���#Ԓ��#Ѥ���NN\���Z���ꔈQ�!.���B~�ck@	�2Q��D�Kz��٥�q��$ *��38-���Tz��o
m'G){�6��c��+o�&��Q�S����	T#�:���f��ߡ��<�:L�i���ɢ/�/��D�����S�������Z�55�u
�~ϯ���L�J7~��^��>����H��>pJ�>B�=@ z�#�U����5P��Ŝ:��7}��.�L���6���{Y֠��6P#��u�B�@hkK#��;���h�h���EJ����e�dև@(��Y^�������:�����3�0�٤��:�Ȏ�M�x@a��0$�.Z��D����'Ͳ��B
0�S"��svv�� �I}�H���ֲ#p5v��	.)>3ƿ�&��.�6ت����ga����A)=0�Ssz�W�*������\�[�ޒ��s����5l{R"�E�N�?�ٰ���5�g25��h���J"�+�P3��)���(v���O��M�׀O�A={q�t� �u���/�Ԕ$�h��9�B�lV
%���9�4.���˕扐�6��&t�zdw�J��q��\O��<+��Ǡ��z9�D8�b�U�E�L��K�+�.����:Z�i��O��U;��t� п8�0Jk�V����Eh�R���x�9��h}R�@�%z��R��`=m���t��X�ؙN�s�尒��:l+���I��H!e��4��I��}f���o:D󖤝�|�9�ZGPs�W�'t����8%��W���%-���M+��'*����]���#U�c��N�����1�b�5ͨV�/����\3��R������Dm��n+VN����d2�TC&�:P7�ݩ�OZ6!~`m"+�\ɨ�C//�s�,�nyf�ɺ!ͷ=�j2f�;	��;M�q��I�ڂ n�U��j��S��]816����`�f���ɦ}~��g}��#�o�5�DM�FJ��r�-�mFi��P+��Y�A��v�`����`k�7YPb.8��e0Rg���z QiJU7�S�i��@��$� 	��77aW.Z-0\9k}��D�m�K�r�温C'f	�]F�t���=��JǖŒWi�G��v:���W�ꂽ�	�p>�îR?�C��h�Ц!�-�Ih�*�o���3�;ƍ�n�5����p�e���7�h���m�Tu_��!ͬy��U&����{�?3����V�5��<�<����S�g���;^Pۂ�M	j������<��&Ȅ����si5�6`�ێ�;!L�d���d|1�8h!�~J)t���-�[N�F*�m݅�ExXV���\R4U�� ��`�̥��^)�c\�� �U�;��M�xL@�޳�kW��u�\ʇ�5
V0��N�����-+��S�k��Rw��f��S��[v������T�*)R傱���в��7��+�$E.td�,�95FBu�9z9�G�̑1ݟR^��oШ��ע14*�O���r@���|�L��N,Bi�4ꛯ}�SZ�WWc���h�$�Q�ܶ�JsA���=�v58Ԙ|�p��ׁ��ѣ�E�N, ��Pad�!;�$���g 
b�+ͬw�%$����C
1�6��t�V#�1x7S��^͌Ӿ��K0:%��b��S0.!	�J�g�y��9ώ&��-�$���H����)�����bn��8C�RΈ�s��z�����O܎��>m�C��N�B@b��:�T5��S1'ԥ���1���U=g�om��-o�>H��?zUpoZ`3��**�� �cd�Oc��-'�Ї��y�9�?6|^I}�m��V�(�7��7�l!?��Z�IIJ���\qիN�L���B���=k�i9Ʀ��A�����3W�{�6f�5���Ʉ}w��p��֋y����� ���o�
�̱D���L��^�U(��+��\�e���=��`�\4�L�zd�1�D
��N4�ј ��t��H4���L@�s(��wb|�j�ĲFj�_ǰ��C�6�q)bxu���8�A��O0�`ާ��*c08�GU�G%ʟ�֧�ʈI<JK�}�Pǣ��ގg!��j�����Z#h��
g�dJs��}+�Xo=�:}�_r&k~磑�p��)�j �&j��L0�~B��D=c�;�<�:;�2]�WE���vt�T�0�U��6Dv�Nt܊V��Vh�.�m$�7�����̢���a�Xy#h�
�5T4�N�k��+g���T�+X��Jv��a��O 5<�t���{��5_Z�RG�?�&:&��\B������v�����
��������6N����w��[n��E�,�^-��m�x;=2|e�i[��Qq��o!�AW<�|�l��N�Z�8��h-�04߁���I^U|��Ae4�IL�1+S�ٮ#�`k�|W�I�s��]�k�>�Fi��K�R�P3)�732��+Ɠj�ת�������e�r���#��D�<�a�Ya���T~�%���a����������4�7�mUȀi��j=����t!�П����������3T��L\�ļ��	��7�����y嶏���4r�7��o�ԩt�w
�Xfk,`\4[�%,bGk�n�d>���R1�V`A:mh�J�)4�]�F����E���N�*���A� 6�(��l���xnԛ�ݺ��߽4�=z�x��.��t1g�PK$�{����Զx�����@��	D����1�9]젶��zm��cؼ���*`EH����%A�ꋹ2�\A������fZ�ꠢ1L�mY˻h�KAx:Z#�A?a�.ᆩ \ �g����Id������9դ�kD��P����� ;���&�uТn��e�l;� �-.��5�T�<E4�"�,T�i/��oZ��U(�a���rz$��]e�|�����w��u��I��7����tB�j"ආ=_wGj�w^_����a���BHX<�>�JǇz��elf�6�?z�|˹m���b`ľ����	n=$�����i=]�2���m�FL}rWQ���p~UP�C����$�� �����楆���@诋f[M~\
-�Lw|�1hq,&�Zr�0��L���qi5�V���v�� ��B/h��|���m�s�x&���;��^�ܞ�:�+;�	g����eQ����IWΦ=9X|�'K��D>lJcx6Y�XAS(O�j��%¾��/���a?l3�X�\��}���酓Mv�؅���˓4%!����K�\��Lx=��*;�����'�蟳�`�3�^��P��3�4�VBι7�6��I=᥯P��G��u7+v�]� '}��L��`t��OJfs�f}� �7�u�6�C��X##^��F���A)CWi��I-xfJ"K�#{�z$h�����F����dE�CMydt=A��3��X�Ӽ�ir�l\Y�;��h���\S�:r�pq7�$��ҵV�]m�p>P0�y�0�@�5��g��8�h"'6+E�2�O��D{koy���s��w�a�?1">���Yؒ���<c
.s�Z�3�H�:�.��@W�m��w�-ŀ I@�7sԑ�/oL����߲FJ��N$���٤����(ÿ��{z���f{��Bj�<�dHt��DȾIC
���uQT��b;yS0��HNT�� �R,՟VhJ,�B~��҂�V>3;����~���re�0�����-ϑ?�+2W���ᛜ�-c؁�4�`�[�QYSu.�����,Gm�$����CG�'h�v<3���ʜ�,Ptڽ?��tю��Nl�SC�
� ���T���Hbr���l��8������S�'~
���m��s��W�}gU�W���}7�ˣ2&�5��<ox�w������hy輔�Yl�2nD.�g̈́�҃=:c��N5po�#nӭ���s�B��2�n�?��ƿj>.�%�'/W�?l��kC���]�~�)�S`���'d�5\t|ny��^s����d���\�q\N}��<C���C?�l�wβ�����q����{�੹4&�h<�����!X\�B*�V�=�erkXG;�,Wr�.9�����X?3�
�c�-U�g�u����9Dy��_�!%�/���v8h/�`��r���q�hX(=�JvNQ�v%����o^N7[^e�wU�[���I�!���V���#��y�R$v����!�ѷH��ʹ҆Z�R�D�n*E?�$�8����������#�l���c��1�6�)i�짯���
%Ll{˝�<лM��q��o��cj�Z��B�-�(Ds�ر7�T�%�H���>G�bf�����m���?{Rl|N�s�"�<Ң@�E�W�#��6*�iNa?��e�$���=����gd��*�?ҘEi6 �}@[���}ۮ��\�E\7�ׁ���$����ߐfR�.X����2���IGYk���'��M�����<+��ˠ(d��u�g��ʀ�W����{_sw�#!c��`�ê�o�/����8ZR�c���p��Tc�K�މ���*M�����y�U64�#hd:Q�ˣ��Ok޴��M� &�*>���M|+LP�/F��Ò{��"�?5���f@�UUZW�/�Gs�a����6��'o�C���d�(�R�������v�h:G�3��`�Y�����<=�uaZ��3�V�O������8��19����v�2I�G�+�w9� �`���.d�u �_Ņ�ei@��k������)!�z��w��菶ߖ<6,��-E�q�˿~}o �>��M�7Q$�盙ձ�����<��y=AS���`���G�N3}���/�V�"$��u�"[o�>�;�����e��f������d/��Ȼ�.��U�|���huj2_������K�i��@��蚜K��*Q0V"TD�	��3z��"�w��(i#Y������8��&��C�`��'���p��m�S��~�)�vA�UCU򻪝��~w����z�:|p�]/����f�l)�5�9�!I�,9!`Zb�C�vժ�8j�&aj+��N������).����X����M�l�D��@iFX�97����m�o�SM�U7�����Q�G���n:���08�m���+5�R�=��}����54�;�Zt����	%�C6�8�%OwY�V_��qE'4ad�=M��sqx�7L"�(	�!���'�(aW���!�����c�����P��Z�$R�9������SZP�&v��Sp��MKzYȷ��:�Փ�Q
e_j"�o7��lϜ����;�_c��i�_:ހ�+���ʲ�/�R�KiW�i'��� .���H��D9%�P�jnVg�s�ߨ� �^��AX����)�j�5�m"b,�仝��e)/ۃ�KK4��*���{ȴ�g�m�����ci�m�o�;���࣬x���s�6t]�{�$jQ�2r�wl#Rv���q����ǭ������΀�����2��v�9����d�M��]OS�ӟ嫦~�k\T��
Ի q�o�Q�!a�E��Wi㪙3�85��]C��S�=Q��/{%A�k��K��"�?F��@����$�N�j=�e�Lݲ���+'���kվ�)�y���7>b�~T\�]�]Rv�E;~���- ������ƵH#]�ߥf�����'MQ ��GL�5�N�Zr��U�,���+C@�Nݜy���7��qlQ� ��G�������Q�T1
�H�c��b�}<B8�΃� "��9D�E����k�q!k�ek������x���N;{hl.����iH����u�M�;�Z2�����n0��������֘Oٮ����d�x�ccnC��^������5��W ��-!��9~��p���/	\g Z@t�()o��´��܂>袷��3̈́@i��"�cQK���z�ן���{Yŧ7sY,���]�?ǰU�tn����cpL�����3� �W	�r:�ǑАz]f�0���D��~�>������*�_����5����+�o�u��`���g���B�;��A�����z��!��Mvet��I%3�Jb�G�D"Pr�O��ē2L��Mm)7Y�����*KluQԫx��Wp�kp��l���]@ܤ�G��	�,�g�]x�j���tLT�m]��\.�qq�)��"����>��`��0���@#aU��h+rG�Fj�g�[|Ac+Z��(bAړ
 P� �4�gD��l��u���cK��ofs߻z�����fH/��<�X5��!�Y��f6<��`������2��'*�vӤ���g�^{v���#�[A 9:C.�Y�I�}�Ț�[g�tL_�O��֡:���C��mJ�d�Hך�F���<'���qӻV�M;�j,W*CZ��zEk��F��૏�_�^{������SN��2f�@M��2�4 aw'�ȩ^�M�2d���$����*-���?K�?�H��`�m��~��eh�+��3�Ce�J(z�[����*9#���N�&�Cc
�� uݒ�)x�εa���4��G��]��0�����p@}IkF�@�:��Kz��O���0���$�1*�X�`R�Y��H(>cM��;.�`Mt��r���� �a_6�)�GJ�D��x��I� ���c��P^G��|K���o��`����1Xq���uG�^*�J:�/vK=z>��(g��2�XHy���jqݶX?{ؑr�y6�C«6N��h���z!��q�sM�v�YR͖�2��0L���G+-����Nt�M N��t`��;���d$�0��_�Hs=��CD�(�Nj;v��Y7k��?6���z�y=��P����` $<��w[x3�s��GN'��+5��Iy��T����[y�Ih�!��o���)�4{��'hPA��Y]�2w.k#�F���qi"�d�+�?k��԰se�9�p/�4��#q_x���7��E@��x][x��S�7��#q��{�����M���(7��wtV`-�Ai�s�;�h�r�[��n����^v�(�֤{/F�#m������Ս��v�7�8(/6�u�-wۉ�t�gԡ,fN�+20��u6A^�9-Z��@�.�5ŎI���."x��ӈ(�Y�h�?�,�E�+���a�KI�06�}��� r�f�[|Tq�Z���@�ߏ^!�/�>;�ÝӁ2#�Ymfs�X���">s�( �ʘN+��y �,]��V���KڬɅZ�YE�L ,���I�I��9���V��[���a�~56����Jm=ڢ���6��2��@�hx�rE����o	� �0�N>��!�h�0ַC�"���cz<���~Cq	&�(i�JLe�774(���졢4ӯ����$��B�,l*iU����S��s�Lҥ����z���[`5�E�d�� :Ll`�Z����ծ�e��6e�	�Vaa��.�WgΔ��Lk�Iyd���-���2�]G���l�1�>�@�F{{���bIXu�G
6ȺQ(��u&���s2Q�e̯��Oz�M��u��@�j&�W�R鈈���	�t��Z؁ʮ1���8U6��5�z|���e
��ϡ���X�C�ʝx(@����6'�m� xu���P�ܣ���˸�R;�,��T���.l��Q�
�D�3�xY��Ѳ���|U���D�=F}/t�U+z�u��&����+a�k{$���v*�yo�	;B�+aM��a��hș#F���MO�ZS�,H,o�}�{�᱾�p�H&bDS�����H�P:6<�"�r�@Ջ�R
��*���q���;KX�� �Ҝx[��\f�u8�ڪ�Lk�1U���;��4v�< ���S�U���8П�Oh���4;DX0`�0;�ڒ��5��#�K�|��xo��A.����F	>�7>_�Ҟ>�8]bU�<x
~�΍���b��g@F�몎=>vK����a�TZ�Iox-�-�1�b��##`g�c�crmU�*_(���~BY�ac0*LtO�TS��pG��[D�����/,2j��E�i+�K��,���i���}8�k�/��+<��VK��ye�=R�D���F}����=��B����)��ެ_e[
��Pm�4����La�ݹ����9G?;pahe�y/6�5�ђozg
p>��eNk_L؊i������`ch򞢾�'�z�z�=;S#��]����p��6�T��|�ۖ��A�`k�����A���q�l�|W�@Q�T1
��ɟ�G����u@��������ਫ਼���&`pJ��;�k��j�&l:7�8`����T!���]�By8с���j�Tt�"�r/)$����g��D��Q$���{[ީ*�ھg�J(:sNB�A�6y5h26&���)����yҐo�Vm�Q�+�W�<�Pf����s�k!��� �D�ݞ\*#Y�������\sڽ�a����)"e��0����j�z¥mLFR(A}}e\�1k�ש�Z���G$�T��[�I3�m&�\���ItGp��%���l�N���aI��vZU�GxǀU�T�P�P�`D��Wx�F���ѧl�S	�al�b��ii ���"�4�w(tF�H"׋��a:�:(2���/�CY�=V�3��y%Ϥaפ-�Jw��.�>��K�St�� k���p���H�Ke��l�/�ˮſ�1圭���A�����7[�g��,������� �	 ���
]��O]+45e�[�s�9[�C~'�[�8�;x8���Q��3���q��Vi)�k�-�ώ��2��H�)H�4$�w�'� ��#�^��+�:	�F'��@��'e�}C����Q3TC\A~%]�5��6]p�W�*l��7mʧ�u�k��o�o7�Ey�����}�N��mɖ�+��!O�ޢ��*�y���;ff�؊�[K@MV��w��t�]me�@7���z��η�G�`���0;dn�O���u��0m�=Z�,!W� ����Cɑ~ŶjT�LR���ea��qvg�����r�B��W5�"���B�MV�\Ht��ٔ�e�4HR�m����v�)ą5�do�uf��k4o������M�d�kF#�p�'euh��Oy�=�6J]t�ǫ)���إ��h��Vj!�1f�_�����h�I�5X��~����LHD��<�!�.078d�+v�1?�����;����x�F�ɘ��Y�HHE8�5��X�~9�^��
V$܇(S�"p���S�0��1cff�-P�4�em�#y|3�w>=C�Bn����<*��� ��.+?E����K�UF�8X���
�E��|t��N�o�6��LA�i��s�����/ n�+����r$��%��Ji:B����б��w �m��>h+Y7�C���B3T�����B�^~[�;)��t��S4�:
v3�q�8��0�5t��Z$��fpd$nb"\�lZI�c��0;��W�Y��x0VX�-�FmJN�tlXh!C9���s��ݛ���D�1B��`+0��S�'���>�n:@
a�z�6����Yum�f#e2Z�'fJZ�xdꄈQy!rëK�\�.8�1���u!�o*��S�z;��e6y|����3���D����E�E�7���(��y�^�h���{��3ٞX�e��������WGw��e?s��tMn��������¬���T3��.x�nI9~-xm)��.��*�� Uc�j �S~R<�g�:)f��Κ�
��'��=��sǨk��<��쳒CJ@X[�Y���y���:fA:��G'�߻�@:) ��y�y1
b��N}� c��j�l�r<�͘iI��)ڶ𬘏I�
+��)��c�X-&��Z���=��|F��1y^^K�Υ�Bה�1^����{�Ӳ��Y\������U�R�2{P��r���=��bn޴���*�&�7�����J���ZP�q����6��i�!�����3�ʷ_��ȯh��h#斑��kP�䣖`��w��?�?T�$K)_�w#1���}&X�&�$_I��}�w��?���L/4y:ȟ��sx޵�3��U�OM�b��&�3��ù����Mʙ���%����^&xa�v�Tw����L���k��mG��6t����G.�"=�
$=D��mFu!�:V�F�J����^�!��{N�f��؈SFi'�tq� �LF�_[�$1�0�%����h�e��e�B��s?0r*X&��~΋�	OJ���b��r�:��a'�`�S1y� ρx�C������nO�I���$)���n����{]Ѓ�k4��&�i�y�&k��*r�ٽt)040:;�?���@lS
6I�*k+�x%��ւz�l��v����M{���r9*4iaB&�n�)�P���Z��&�N��)���) �8`�b�=��-P���l6�1���Y��D0���$�s/�Z65X��c�i�;~�N��=-R^zhfHLv�X�5>(i;�H V饺��.T�!8ޅJ2\ 畬�zk�FH����M�$�e�1萦s�7v���S�JC��jg��EϦA�,�Y�F���lKG��I>"H�Yț?Ah ?�g�lU��a.�!����k��3�k�f�"q�w6H1E����3��淮�D�<�J��Շ$���w}����]>�������!�o���tb�1yZ�/��33��=3>�a[��}�i�b���3�d�N}n٭ΉYW�0��0�g"!G�]R,��g���uv��'�u+x�FV�'D_�mf'I�_c�s�>�xK�՟;�l�G���ݒवT(e�bM�-�y�����RjG�k�n�~����nz���/+W��)��������7Y�>T�� �G�����Q��&�t[�E�vT:�7������[�,l5GX.v��W-E�����yN�)�HH󍥓�$l�?�ֳ�(���>�Bx��r��M� ��O��:��
	r�C��q>�U����ԕO	,g��5�T���k+��H'a}�wy��
�����eX�������񸕻ap�S���ɗxR�F��C6�Ak@������8��[���!��̨�.u�j��ڬ1~����7L��C�W7c*��d>�	-G����oH�d��>u	p�[�ވ,�.��AY�w��p|��Jn�_�T�ܮYԨk��=��G��=�lO��D��}���`���(#�Ϲ�H�Ro^�ϾJ�^�w��0���̜�h1	�9C5���DRe�h^�5�)��{��	>rk��p(ё���2���\e!��VΩ��To:��V&���@1�_��ݓM�����������6��S�����+�^���X7R�#%�g��3�d��>� !ث�+��A�tD%�yb�WY�tA��@����@�d1T=ٍ�$,�F��f(�n.^�R�R۬���[vC������ɲ��Q�8�*՗6(�	V��/��Ux&�e_b�Y��*�a�ϴ��X�φ�#�����b$�?��fO��������ZD4y$.��i�>���j��'���;Lk��^<,}�]��]+�}Mv1Cag&�u�Ԝ��F�\OS��~�X3��d���8�����,	 A9��8�8SK�����斦a�ҧ{��tW�6�H��p����",\kH�������oC�J���6&ɮ��-��G >q���T�p�[S�pܶ��0�z�q[��g�k���9tzt�^#?����ܾd� Q�� o��3Mj�1��B3:�z�|H����<m
TP$����nԻ�`f��g^��{(c�C��7y��(������E����f|�ͽ��9�	����s�Y� �0{���A`��?� b*�;:<�����RB������!<�2���^G��Q(�b�����e�'p�Xvf�r��\ɻD��֡Ѳ�st۝>��Tc+����P\Nn������ȓ�jN+����,���Ԃ	�3�7]b�Zظ q��G�z���3�g�'�u/c�>WY�x?�����i�)� K�p5���-냔�R�mW�**ӻ{ e �:���<��� ����W���{��swn�n�U=j�������\'6Z"�������yz�&�Џ+�˰ަ.�� ��I6Y�Qs��<�X@!:��/�J�ߢ���=�<�A�r�f˼�F^;2�����^��;S(��T�ޘ6�I�����Lz��\Kz��c�:6'$�"E�Boe�w����Ӽ�z
a�P]o
|l�З
���O� ��F�T|����;?[��[�j>x�����|�EId@y 9��D�HK߮w�D�0B
�l�lȋ�����?��wj�'޿�x#`�[E���.�����y�����C��V��wvK�I�X{��^Ug��R�C菗�,{~/ts�:�3R��0:�,3^�_;�\<��K�y�I �,�I���F	T��6�̀�i���?��N{j#�T�P�����D�e��ĝ�{MȂ�P��,Dd���8�s�B��[_d��}�AF<d���%�)��%��?��:�e�-u�[��2&9[������?Ӓ�@[U j�O���	v�N)!��x$;#@�w��TZ�\���)ë<_��v��s���0�v˵�d�~P���w�^�<+xr��{��mV���mЫ�|�$Ѕ� ��g�"S��|��$���c�+G'pb\j���
���fh�)����Ps�c�g�z#\�Bs���Q��8���x�VSM&�ø�H+�.1�.m�-�&W=�g�s�:��5��[}�ӈ��nߠb1�D��:���M�(�	'b��ƪ��8
}z�|��uI��aU+�c�ej�&._����SI�)��:��0�(Xm�s����-�]�e4U!�J�gĶ���o��W�B����+:o�D��d^K�	s �_�G�K�<�͖tU�@���D����{wIh�wu8Fz���[ ?XG���v���;��&�ˍ�M7׋����h/ת�I�0�}�In��r��L� 1��G^���v��E��
O�h� �w\�e�)'��w��ڧv�|:�m>�i�x���XR>pͅM��z�;{.��ys�O����	�J��ok��~ h���8Y��>F_�5v��,��khE����9"ơ	���v�+Л��|{$UQM5G��q�.����,��F���-,�sg��������].S�����E��X����gu5z'��b�@�_rF����K���L{�8�*�E��l���6sr��I��5���Nyl^\�&���L8��q��"�C�� :Dl������a���L�E�&�{C�7+8���DA��I��y]�g�oK1ΚJm��q�i�J��pQ?���+Ӭ�x�/8����]�/oEhK�[��E<asH�3q�a���a�!��w֙*�O2���
��g��:��6)���p,z��R����1V��v���η��JV��̡k|b������)4�?�k��=Rk��ɡ2�O����A�"��骽@���,[>��r�g�����#�E�DjZ�jo�E��%F�\�~+�ƌ&~��x���~�BUn� o�?��Cϸ,Ӑ�>�f��w���	ql:U�$)M~�9�}~�K�yEOB���>D��?��a"{��u&ZK���;�ґK�&�1�\G��V
W�U��g��B�D(}���N:�nM2��u�lm��w`w��-N7���3k! P���HI����G���4^{[���]n[�՝w�ɥ�_D��8]��,)Jĭ��z��O��{ɱ�~���:F��ͽ�j��G��N�,!݃��.i�%S[�/L]2��\�_^,H�h���~��<�{��Y:�}2,��@��eʚ�\�B�F����<dERWa�aG��!`%Z�m�Ḷ|�0bn=���f^`�_�7�+��Eˠ�7�T��@$.%��s���w~E��v��aj�[�1L�h��S�7"�rbh��=��ro����;�����~��T[dZ����R���U�qL]�hw}�h�cR�{`N+��hR���z���Q�[V���3&���ڈ��H�}οy��t{��ދQ�3TX��p�sf>K��$��P�fL_0~L�hl($|$z�S�3li���	��F�#�I�{7�&-�D��a:�\-�Zn�B��ő�k�ā�S�+��v�]==�~�[GA3��}�di��d��n*T>��We�>�|B6e	ʡ��a�p��+�ޕ��+���L��«�c;	�)[��q��R�2��y�.bȄ�P��@��Adn7`;����`���q���ݱ������gK�5_�\#�Eog�W��̕��
�$5"{�����.'��N'���m���R�^���������/�ٴHo�e�{�(H���W��3��'��/H�7��7�լS��s����W�h�F��D��I����Ǳ���}e�R��l�x�t"z����tB`����fnxQ_��R�Ʉ$-w+g��N����A$��#�&���c�<d]{�S%��_��+�t�$��f�Y6�/�iZo
K���!����avv޻��C���G���#�O�/�Kd�`�i;C�>��q��).l���Jv�q�z2���U���6͖�q3<�F�Z�����s:�h�K����C��r&G�ax����E|j��?MV���#ĳ�w�"�l:յ���t��	ɚ�b���9d?��z����Z�'�K��5�5	yW��>%��Ԕ��w���9�.S��WϞi�c~����u�W�E����MS���`V���S�:��=��^�z0^��]���V�n���B�5��Z;L(��`�O�i���d&��jI~ 
����\e�0._�Y�d�If�i�͸�蘊�ץi�G����8Q^��^�u㽤����s?���s��s�ݨj�"�W@C�?*h�P���)��M����J���?q��/ɟ��3T�������|����&b�|���nВHz'S�c"ɭ�B��N���2��R����(n����N�E�/�3�Iv]?P ,)�xt��Ǒ��k�e�G+nnq��5929S	����=:�� /|:Nt�ʮ���}�	D���8i/���X+S}�^������r%'�-���l|M�=D�'���l�<K�߾�dE���b1�����XE:�w�N[��$y��=.#?�q���<k�k,��s�ʮ'`1�w��Y��p��ֹ(����{E�.���	�Z���^w�ᦿ��g�*�HY���ޢ#eYXA�ge�=��b��x�˼���6�����Ǆ�ըo���Fǹ�_�f����ba�ѷ��]�xV'V��l0�|.R�5	�����t�+xBb�G_�����*b�7�oq���ޖL\^�4x��-i�G�I����K#]��0�q�`s2-B�_�:�Y]�����ǟ�0�@!u�Ѕz
��+���,�����^h�NX�4�{Lnr{BT�c�e���v�1OII�B�_pR
]���x����y��5��'��R��p^��h�vq@ST��X�k�5�v�p(�z43�lQ�����J�ï�!�[�}�m��r�@1d0�9Ƨ{�zFq����).Ƙ�F���Δ� ��~!��Ԍ�7� H>*ё\L���sy��m��*�s�"��y�p�wT�Y�d�a�R�c%�Mt	W�����2��.�����l1}������:�x>SH��ZQW�ơ��E��\6�HC�cէ�6�0Ӡ�S�mM�&�J���ҵ�����V/7xY�"��N#��[%R���{�o�����5K�5���c���(!D`��$V���������s����l�'6����E�,��$vï���B��k���ڻ���~j�y,�%�ƚM���7�#i}4��|��Sw�8�9�6�:�
�d�����P��f�2�hL�~+\��a��¾Yw����|��<��^����2�9^���c�������I_|L'@U�'�jU����ʤ���Cb��$�/�n}�',aε���8k�uZ<CI��"%>ȡ�n��y%ݧ&i�J�\c�b]����C�XGH%��X5�z1��<kOi�+�¾���>��앐�p�V�v�`X�9×�v��8|%�3�  �u��
�D�'G���g�c=�R���F�p�+���Wt��	^u�?&s�MP��P7�n�-^�������"Y��{�>�����#{vid)�53���J�_IW*��-d{Xy�7�Iyʜ$��sV���%Q��K��4�[�qsXD8b���܆z5���uw[�3i͌��� !
2`���o*�}r�C;͸�'��> ͔xdC�æ|/�ב��-�Iq[�j�H�=��xlof�U��BRY�}�¦��E�M�Q9,��F۞k�yV��������Z$����U%��\A�P�M�Ȳ���D|�����w��0��!޻D9i7z�C��X�U�x� �f�t�J�w�c�A�����Y��)
k$�B�6*�Ψ���e�8&=. �Ir9���m�:A���
c("��H���L�73����LKρ��q�c�#*l���-����l���_L�,�����˯:}����#��u��6#55�{8N��+w��B9a�
��c�bDr9}7K��"1�Q�-��A�tX�;�p_\�k�'��Z���יj>�{����i���֣`���-,1I ����J��\���B��p|3"����nU�1:����6��_��/%���q�#����Y�� �����Z��Q�em}�uN�|ۓ�˔e��	X7�5�>}� 3�,`K0��2i�4 o*GV� �/5��{ĺ��������}��v�7��?��U��D��(�J�͛���w,MP[�Pg`Z���r�]0��\�ڈ�ȯ��5��2#�7ޛ
*��C����Rl�ʇצ��:���cw���t[����D�S��c���$���R��J��Q`�î�M��ch��2$��8���r�x�~��%������K(�?���N��{8o�:OTlg�KQ�ї��zbߞAE�iK->��G��R�U�Qc�!�"����_���:8D��v�AJlN�+FH�Qk�v[�(J�R���Ku`b/+c͌���ڃ�+ٺ�W��]n��-,l�؀�ʏ|v��;�~#�I���������-��)cI�mL]��ݬ���Dt;� ��߀��E����h$�\<��m�_E�4���-���IвFhR	[���d]���܁��d�1�r�:�jL�B�:�⣶ X��?72��f�%�?s*�MXb�-�-�;��)&��*͙��z!w�h�=��W��CT���m�fNT��u���P*�&�69��`*���Hl��¥x���w��	wu^�� �mo�X'�_��,��S���h���5G���ƽ�@2d+��.��Hϟd�Q�B^�;}o���>�d@��� ��nf�KĦ(��Q"�����2J��+�94_� R�9��� �����*�v#}ˮ1^���P��m�&/'��lLɁӞx��k��ş���1f�v����N�
�F��m}�"�W��Ѷ�,Թ��|��jQc�mv\���h^��V�x��sJ8���m��ٚg-6�::�AzwL�h�%�n\̖�h��� =���;�J�^k`�o�m��N��bc���٥�Wv��|9t�b3_���fG-F͜Gs�����^�;��߬{%�)�xY8�Ȣ���nW*��� �l���A�>sX)��\;	�����Kd|�WJ��I\�O|��80�F�Bg��F+��9j�lÕ��f��� A���{�<�E��R�s�>P�f��ad/������~���b 
9� ������z1��M�ǒ�b��ߤo�3�f��Y�XWc|���-��� ��ك�i�|�t��n�H�`,cu����
� ��64�
Rz������6xU�2�"�+�V瓛���Xaw�:�����(�@�폨�D�,=?E�cyǯ{��]�cI����3Yt�X!�ҭ��8zw����!�=j�/�@(�t�R��+{��b��f;�ȍ&p�Pm8�Q)L��s����2� ��*��v#;�W�~�x�\ ĸ���G�B��Dr�w��:���"���ص��A�%�>V��6!�
�t�>)V�.�;�F��1��e7���}�����K6О�gǞ���l�g��-�@����jnu-�bS����������6/�2���N���Wh�H�mo�l�,�H>%e���c�sRP�A�	����2����	j��v�'��W��>,��%+��וo=��9�O�5��9^�!��_&$��v�a�P���Y�ֳ]�$;B��y�����̗l�e�ȱ�i+Rq�px�����j����.x�,'�@��'W���c���qgY�8���Lf�ߍDկۘ���S�"��>�uNvvOa}5ʮ"��]�O��s�M���W��6���nm�y[F,�SJ�oV�S�Y�y�$���qvAIc�y�f�1a �|e %'S|����(pJ�a9��+��ٮ�8�4jAU��5�~^�:������M}��V�0���!x�2b~�D��G͟U��2'�t���GU�C��]Fdw�3��@�K!�����,��$�M��h=i7��ƌ¢�dN�|�NS�RM�>���d!o�g�Pa�0���ǲFJ�'6�<��s���[�2ףfCC��Sp��uu��!4@�3=Qm�[���j�3��MN
���\�׼��s��8>d5*r-!SZ Lnmi��\�*��|Z]����V�{"�ɀ�U�;�(Hp��������G?��C���Ď7�6Z!KD�q·u��!`O�ѧH�r�n�U����=i�JAL%qi�>��9R!�(����Xp��F�j3�z״���{9n�f�msD p��X!�s���Y��|Ex1���<靈*B��?Fb�(��>5Rp�˼�^a�X���T�H�&OZ=8�U�#*�/��K��L���e�'�cǛ���HVZ�ڦ`j<��v� d�i�+�tK~4h��O����'�_�p�!L^�]Cj�:Ar2߀��s��j8��It�X�e���{Ow��m@�Ҟ�S5�����H�Oe����H8{���j=�U5��
8tO�����#��(�ޜ�Q]/)��0uoQP1I��ʤ���pk�*#�-M%DN��ee�:�����T��B���߷�&���午��E�g�������#���'�^֔8�@�9(a���e�Dn�<��\Ro�JA�_�����h�a<��~t�'��7���x�;A��D&`4�Ә��h«�fN�1�7a�j�q+������4?�E3ڑl�Н�>{�y`ӱ���X>�-ַk���#��ǁ�G�~�Ћ�{�\݋��5�D<�d�<JibO��0����*�!Źԓ�Ҧ����)tүѤ�?坸 �4�f�N�S��b�4�.!'�����}ۚ���|>e?[�͑�ȚX~�!���	�l�,���K���+�ToN�G��/���IE�SAr>�Z�0�[?����+�o]]W�������>0�R-�k���*ҁz�bR�$�*�oz,o���k�^�yd��0��B.��0;zO<!&���L �����*�f��}̽G"Mf5T�-��)�\+u&�?��o6�.��<�~�q� ���h{�E������^sY=�H��wTy�meU.���U��	�r�H3����8vrM��4�	�`�0D4���!.���f{�>��Q�=ėy�.)�D��*��s��)a�1�_!���LũՊS�:\��>��;��ݸ���C=��k �-=�i��,��_�>�A�|�l�����<���8b����������y஦�6��Ğ�~�S� ;��t2��=�����|3�U���͸k]���'�F�X;��p�f�~XQ���K��T���-S!���>	�Q�?�`bhx�lhS#!.�­Ǫ��S�3�3|�9�]c��_�w(W3b`ww��r#��@-��_1Jd�Y��|���H�JI�A/ci!��8�g�,3����Tc�g#�bD��Z5�E�����((b�H���X[��=
цVJ��/�1hmN�dĉa�0����4�s��?5�h��Z���5���4M��v�e�=+GD��:!3��'̡D�*@�V}>e�����F9���ՓS���}.���
E�A��<����ݍ ��:�;q�U�X�*z��S���ƿ$�c7�e�3�KY��Z�����}
`OSx1�h7�P@��tl{�>7ol�\�̋}�yJ-�WtZ�y���t0w�i.��|���Y$$J'���Ks��
6G����ז-JU:�QaN2�#�s�' ���'A���-�u�&Wd-���2�G�	�����^��'?��Am!B��Q����ķ�mpV4Hͺt���y4��}&;�iL��N鐃��J%�����5s��G�q�u�xX��:o��D�y��k��Y�wXt4I�����s�ƭxC%Pl�A��B곤Rs{_��jG��a�L�s�7S�0[���)�z%�fAI����s��®h�����Nb��V��g���u�PA�RK����mU�t�l�q�O���u_s�2�Nֿ~�3�?�Be0ևQ�2&W��]~�V�O�oz��7� 	8���ۺ��w��j���A�h#��'�������U�ȫ(Ȣ�Uj�����MG�]�0[(˛{u�1H��Y�;P�{
Y5�Σ&��=?E�D9�P�s��m&c��NcQ*�q�h�0��c�JM0�a��2*�>ϋ;^ɂQBH�(ӳ��C����l�w�1]�-f�Q�D6FY��QJ��y�TbI_QBƋ�	��ʗ��M꿨/+� �!��!P�T��C]�~��M��f���h]����2\�]=�e�{�s�w?DX�W?
��y��?u`P�e����ʉ�����������G�bd�2b�U����ծ�
"9��X.�����0�����*�̜�T�}3����?�%�`�]U�����p���:Lo�-u���ʪy?�P�����������=o����#pq��Uq�Н:�֮r�5���f�`N 0��I/d �G��t��� 5g1���`�g���H��6{c;e��4� ���g������i��g P�-����)����b��=�"��D�^�⃤��bg��Ϙ��z��U'q��^��MN�U��ڪHt�Me���{�,)�8d
)��o��`=H��v!�
���A��ujۀu\+ �:�:������jZZ����W�^�I�\��T9f�K>R�ήN�Q�3���ڴB���0�}���t�:�
eԫۥ�
>䎨x&:ۿ�� S�K������DP��bpߠ�m��x�#��L>3x9i@p._�],�=�z���q`�~C�����(��������7���$DV�{�A����a���O4-�4�y;��i6H�D�1}��ӸǴ�'���D4�� XU�ܡL}8��W�ǨB��Z�K�+w�u�f>����y�ԙ�j�< E�{T�xZQz�����Df��6�Ή|7#��K�)@Է;)>�m�o`j(U���q����<��pdtL9�R//&�@���u�(��eP�"��!�Pg.X�+�xϤ|�ϠI��o�����gT����SK���ޝ4��עt�|)�����&}�>j�n�����F�)v��Q8���H�]����\�f���?p��'aL#�N��H��%}݈�V�a��H]cF�p�қ�q��|���]E_굁�����;p���` H0U���Koa�-A����g'�Ԩ�4�X��В��䴳ǌ��
(��F=�NC� =�dU�M��G�m�ڪ��Y��ir���ٰ-�<OK��3#�c5�E�Ic���@?�o�+�?�F=�8��\5�#qԳCɸP��Kf�4�#d����6��K��k:�7P�[�G,�[��`��\[�~��B!���h��Z���nV��<򝕗��<0i@����cw��~��[���9��TQ������d�	���pۄ�h���aG�}X�Ψ���M����0��O2q��k�Ӓ^y�!���n���0O��^���	���_��9k��l�����	���1�uM1��%	ӷ1�e�ʟ�����~Dxi� }����y��݅�)�ҏ�Y��s��9e�xL�����"����EpǨ&VL#:��%�*.�+̽y��%��'Ôe4ݧ����9 �~_bI����1�G"T"J<2\;��"�jl,�dO �O��c�b�]�o.Bo�6��s�/88VX�U�5�i���
x�1���l5ބ�FD��h2�U�^��|�V?�S�T9b�>�kxU��������w�1�
{���� 
į�|��v\�w).:�B
��x����A֑���	@x���|`���8��?f���n��
��5�^#ʊp{՗?t.�$\�'  H��3�I)������uݜLsA �!�OgAv���Ԓ�>:�����94�34���G~��@*\�mA�`2̋>��%�jZ��|IF�J��%%�0kc4��c1G�-+5�P��NVt�)���j��i=p掐m�f�|�&���j�B��*$g���f��/��#d}H�`�=P$ȰD�a�䴔���:���-�)����=���h�7����`��� �]l`����P�<eK]����M�iU�U0��Rʦ��<k���78�Ef#�X�v8�b����u����.����?�&n����m�1 ��_Af�<:�X��XV��� ��7�^8� ����-�L�M�#�ܚ��q�[[E^���;GDiTڻ��1���MR��O]��A&8��L�{м���~>�_@�8"�=��F�Tq<�8���d�c7<il�Z���8�[���ܪ>�P_�p����?���0��d��	�p��}v<h� �bt�������	��v���Sl]��n�O��3ݤ�G�(��d{��j[���E�$"uz����o��A�HIo�Ur�t�y��=�(��n@����
�f
��X٦z���`#L��ݟ����Ϫw��&��B޶"����ֱ��Gh�a`�?�������s!�F'��U�b�-�����0蠅�Y	�C$Y&'0�i{���&�o��a�����w�kZ����87'�v�ƍ���x�c����`M�&E�W�6�fJ���2��l��ru Xdö���Gb�l�w��q�u�܊�����.ĐL�4χ����s@�1"v��Ԗ9w���?øHl�B��F�z�q���Ltŝ�&�'<�	�jeJŧ�����`+����;�M���@��$z-^�s�V&�m:��ΖK-�r%��m�BK����\ �J6���u�)�������z*jvO�R~Eט2�W���Xg{{q��aP8�혠�ώ���fהw܁JCR q����b��H�3�Y�5�2lUL\��1����ا�����a���-7at�����V��Dy�&
�1�7�_���t'���5��Fgh��#��k9,�w��N��@^��ʘ�L�J�9A������̮�!���=<��ȟkk��4G{&HS"�ܒr��4*���m�{�/˼����lºK�3W�0_��lY�M1�`"n��Hx���|�dX�,$?�+�'פ����th4�I��=H5������RC�>�}v����H�ɚ�(�E�o�����g���r��|1��.F�w�T�r�n9�n!�I���%�|\o@�k~��x�^����suXJ��Y���h�I-�PGL+i��R�ΝRcɩ�=79B,w5<�s��J�H�a�7��IO��	�'�Ə��H��#��d6@�ܞ�J��`�KS� :���s�L�U9�N+����J['���$G�j|���5��
x�oPg���y�)�
��NA�>���Z����>s��=����ҟ�ġΥ���-���4⩁^��U`gԆ�[l0�А�8��>
N�ŠZ�!�O�>P����T�s�4]�-#������|d��Il�=���E1.�c2�Rh>2��Da�V�-�}�D��I�ZKN��]�E\H��OC}w��B��zpw�\5��:���nCfT�J?�];���l�~��b�Ny�^IU@tX���7H2�N�;lM|�^֓�v����%��F!a�E�;Cd�O<�B�����-@��n�G��!S�& n'�]�[^�7�q_y|�$ �%:K���A�!܉GV�-�x`�?�������(H�I�h��/�ݵ��@����zĮ_��N3�j���v��T�A�@�/�i8��f^�ִzC�a�N�����4�q���p-%��G,�D�jB�0i��f��}�"���0!h�h�h}IMڵEDB���pfKx��YX�C9���ќ��o�K~�G��Pt�vK�B�,�þ�_�R����v���6�7S�w
AB�<y厓�
kL~1QR"���������J���P�e�Ԣ��Nk�����!]|~��>T\i�U��Z@b�����<��vD�%G�hʯXc�ػ��m��'�u~R�us�EU��/%�'S�e����<�%�qT��)��#�I�cɷ7��NT���}a�H��/�E��">'X3�\�rN�� Ql9 �JF�R`'!���@��Tv,�<n�j��(�d�3��}����Պz�P���WZ.
]O����s�c̊�vd�3m)ܙ�S�	I���>6`^#�5��Z��=#`�|@���q��0E��pu��<�P�q0ji�ޤ�39�6����j�oՠ��/��J�`�P��Ϻ]�-��Q���2�-.�D��� +�Z�R�t�}(���JU �>�Ս2hk�h���El��a����_�%�F��SK�s}�a����E��S<�u�� ���1�Qڄ�E�M
��*�y�R�8�/�.\B�G`
�K��E�@X�T�a���0*B�i�q�_&����h7}���.\�# �S�Ȁ�|W҃Zw�LW��ȠV9��!'�IY�{�^} ����M��O���uuΈh4U�@�B�9.�Z�y���Zi�lȇ��]�-U�B]�e���'�+�e�zQ&Z�_\G�:�E)��T�߭Zz�>��ܬ�bT ������=[��������� �)J�^���c�Ԓ�8\^��.�֗]���1��:���p�ٟ^	�.r�R�x���Ohm�7ϋ�s2�t�^;tD��'�?�:�A��n��+�x�r���1w$�77q�QŊ����\��?�4�-��4��u�v'6�@���O���{Η��5.�("Y��8�%4p�\w�Hz7�*F�]-kM�}Ka$z�Em1����OK��W
�EԙCB�P�7ݚfV���������=��G����,�KU��*in��HЉ�&�N'�$O!{�J/�l$�_v�ifZ&W�o���l�(����].#/�ed��\\��I[�����n�ȈG*�� %�f�-�X}�Mo;$ؼ0wok<A~����L�kjWVJs�Q���w&O�k���8(Aa �Xo�D3� �K9 ����[v��v��j>�� �-.������͇�q��LWV
&rg�G,P�5˗����� =[�h�%̈�2=|�Ѣ@�������.!��Fϧ�d�j��� oݘ�-^O�s������U>*)v^�O����>��s��j�z�w��e�\��用.NF�T�x�$��b��y��:3�͜�$�R� 4d�0�#�K�Eك��&�@חF+��9�1�74��#z���"n��aPAT����9a�����@�QG�^u%:h4�ǦE �d�&�u�НY�0M�)�ċB��*��"$ל0�_DzRd�sp���ҍ�������qF�3l�Q�~HL/Z�V@���]B��fyikV.(m�R5���Z#g
���.\`?ݚ,���Pyf�2)iH����A�'���u��n�"
j�U�νhNi����x�Ds��
FQ�X�`D>+����˨���fV�}M�
�ʺ�׫U�VHI���o���M��3��w\���o%Z}&R�xx��(�V��Q�`���?b�YB�&�'Y���^B�.qjM}�ۑ~v��L�6,*e7���gk��D��:�G�XР20a�_r����\!	����p�<�)�j2ߑ4=�*]·FS}�Y������گ~��z���vxď���S.G�M&���̟#�@ vN%%����F�l{]��@e��������b��������z��������4w��5�	��G���O��ee�B�%��[q��B�%T�����l��{��L��g�'-Ɋ�`�&	u���"5�-��N{N�J�%/�G��L����8:�u<2S���?�;	�����w���D��($A�/��I{f�S�� ��S)�־���-�m����߄6�}c����J�6���@���{gEB7�װ�������)��5��R'��z|2���tmh�o�``+���~��]��Rw�"�z���c�s�],���_�X����g�~�'�F7��엡���&�\�9�˛��Z�)��X��.Χ%T!=�i���Z��Ӊ�%t}@�S�K+fζ������L0S�����(��_!ōM����=gDeȾ^��!9����, �3%���#<�omf�
 �v[�l�&���[���m��-���Ĺ{�T�{_�ND����έ!�V��3_U��u�N��onW~��C&�@�]��j��J�+���Z uZ�ؼ��C�E��$N^&��*�y���Q�i�L����&��9����>�2[���Ơ�x�R��M58N~��/��Ԝ�l�2�I����ct,텪����O�ډ�.��y�4�Z�^��q��/|������Q)DE�7X+Ȅ�]]̈��\R�b�d���<�&0`��Z.��X&�}���,�c��QM�n�� X_��o�=1��ZU��Fe�L�C9T���"=������%�7��Bl`~���b�����]rh�r�ɗ�c��r�(6 ?���;�`o�eP�y!]ES�~v�Q���?[_�*޻zQ*&d���f����n`Ϡ��E�d����3��
�ƶ�\'�b�}�}@1h�^K~nW�aã��K+���%�WF�w&��G*0�_��/g��hHU�d�����UG�������D���D�He#���?Im铂����ΐ����7�
KեrJ�纋�T�$�P������o�nIM�L������7��I;ɼ&��p�4�+�.��k}���(H�Pb̆�@�y�.�9
(��c�.����L�0�3̥�	�M����P�G��;�(NJ��6���`�З�j�j�r�x�캖�{ρI�hE'$xR��}Y��*��d�a� ��n�l,��z:�~����2\���66�Z`�3��c^��[�n���h���� Y�E,�'�Uعq��Wc��>�X0++�KE�A��~�[��wvA�=����]j��K�B���	��'b����Z�kL�f�6#��{%�KX�f���C i��T��������QF��ÏY��P��A��R�f�U4��" }��{����ib��.�n�k�Y{rJ=�Z� ډ*0�<����S�f������f^K����i������/�KI�.�-�9l4F~.�[Jm�^��^y*�3U�(�^G�H��o��\&x���w���� hJ�O��'��d�G����7ڷw�i3A��z���$m�Z��"�u�Z��B��T��<��Uy��R���yU����.�Q�;�D;6��7җ��,��È��Ĺ*"��p`}`�"[v�����]R.�{�d���k���Զ*�9�+i~�-	�Ri[��B,<�֏z����l·��'��X��E֟u����N_5gu��u�q�I��g�C��RA��o���g G����u+�/�}��)$�>l'�=���>8Cj4`!�+<�^���M��C�ҋ����O"��fF�r�G$lw�ֶᛊ����u�Aڠ3=���s��t��"&�ۗ�S�u��Z�Ɖ��Dö��a�s��K.��/eڂH��:YA��#�����K��I��!�Z��F��s��|z5�#��p^���6��4u���}X��|r�elM��I�ҠQ˚:Z��Η��x����(<+��(Q�`-Ɠ�kv�5��'s&��ߕ���{ӂ��G���ק�.6�:cl_�%£ᐏ�%^�?��/ \R7x�����_M�sި��⻹hNw���ۚ&\���yІ��#�c�Z���(3���mR!�c3��T�*��v`?�//��������W�c��2r��:���F�@h�A�_'���-���p�^��9�n�TF�݇��4���u
Ҷ�rq���/]n�w10�*r�~vQ_~��'L`��+Re>�z_T�JnYV�[��:�nbd@��%'�Hȱ9ڰ�mL ��%�W�n]�-F��Sx�F��V��>��Χ���@���4.�_mi���(�A�jvD����PוϮ��}��3��Kn���~���pI��`��YRr�㆖�y��M�窕L�]S���+ݡ�un�sSitr�t!v�Җ0s�(��_��J{I�o����<tl��C܃9Q�B�\��ޢ4�%Lx�����'��BIn��:���8<eC���>,�j2�֔��0釯M���Iv��2�MʛĚg�[��b��_TX�t����o�^Ɓ�p��JX<��]K,!���i�ǃF�M9E���`��B�I=�2�Q��p-� ΁�k4&�
��V�2B�PI�����D,?�,a����F���ݞ�x}U[�)y�-0�ז��e���Y��ȁ�~��?�}� -xX��Y�s���H��W�g�u}Z���>b�f����}�������J�'�0�n��Ƞ��e�������~&x*-��T��95k�T�ӝ}0-$qT@d�?�1O\����j"6�g�vRj�զ, ®���Yp�9d�8+k��7�b�w.�Ϝ��8�G��P��O��^�Լ���8��1�2}���gi�TXz)X�/O�֣j�f�5�v�4[>� ��-F�p���:i���ճ��7�����
am�����9���9|�t�<��|�p����@x�ә{��o�W�9t]��h��e��*�b F(��9�]�z] l�8�	��%%�U+j�i�I ����W˷J[�����cZ�7~$ӗ�����03������j��(GƬ�!��a�����{�.�7qJ-9�U.)�{y�G͂-r ����+4p�!��a2r��=��C�?����T��ɫ����QH&���r�jU��ܿ�!	��Ц�9��)�>Txq��l��E���?�	�L���dyy<R�bmv:�*ÕX}��,���9��&��_~W���5|�$�,K��I#3
�X��ef�5&���N��� �!��J�.H:'I�q���WkH�2B7m��J�ر��͡d�tʞl��=��{����BfT5�>��}x�A�%���Q�/ԙ���e�c���SV����&C� �(��%�&��l�Ǉ^h!�	:��\�ۻ/"����QO�/Y�I)���]�q����3oh9��z�Ƨ�A��{^b��x�Fq��ĈG�.[���:qL��~�<k���a��ߕ��҃�r�Q�^'�:վ�G$�D(�eZW�F��t�2���(���6{�ă�liӛ����f{�V��,A�ŏe�c�䏎H`.w7�>аi}e2�wE��)�i<GW��?����}V����N�ώRB�,È���fM� �eW%�*��>���8��2p��0�\�>���7�[�����o;��)�n�b��m@��}9�m#���,?1*[j��v�����|x�E�+���Ny[��z��hӊS�sl��|��48<�r?'?�!�&B��o��'��5�&��s��Ƈ�E�M�O)��C>�M4��q3އ�2O%-�V�О"��~���ߡk�B�B�@).2�T��#�X��/���2��y��	XV���8��I_�lY�%���MiQ�>ø^v]��!�ÅpM6^X��C���6���{\�i�}8�d��4�_4���vf����7�!�r���wo�R�TʴGdIU6y��^3�A�';���{:8v��ԏ�u�d�<�N�s���3�F=W*�C�����:�@��	H
����'�7m���:%�R�Ț�&�~�7mI� ��W���U�:e^�\�?A;�n>���dB�X����w};%\���{�l������3�����Xh��?��K������Jr�\�0!�4iT\�5L����Y��&+��|j<ʞSGv��?�� �C�V=��o��3�콅ܥihn6!�֖����U@ �л�;��FX�gQ+���b��3�T}~�9y�,��e�_���n�ǽPG_���NuB� �����U2��|�-w�g����]�w ��TR��������:�'��"=�x~�
���f�(��{�d?;�g-����O�Ekx���d�l�Gt�������\v��"=�s�;j�d�;q�zܤ���"д�C;̙�3�P�I�R� �&kP�c��l�=�ް��<����?®��l��n���Z.����9�Q��|@(2,R0���j���y!�HWq�hQ�ݵ9Ŀ�/#�ȉ}ٶ���݈E
��o��]Mm�Uf�	����7~@��,�j��v��F���Q�KH����9�R�'j���P����4 �$�b�kA
?��}�@���O��v�`�x~���v��fT�?����z�I>�=St�Q7'��������L� 2H�~j�^|���V�H���Q�|����j����I�QWm�=ֵ���k��[���~7$W�^dי��(O,��l?o/�V +�]x�)~(��B��j7�U�4�if�[���|���#%(� �Dr����1|�r�o����� �/w8�?g�1<{n�o^���K�~�"�qi���Pt��B��&*��D����[���|����]�uM��㐎��p�N�ܚ��'�$�yŏ�����2�^�K�Gr D��y0k�^B������>������l��/Π(�K��.�+���.�̦�o����	��Il�?y��x�!��	dA����T�B	y��B���k�� �*�c��L+iQ�+����!KV3�e���I.\B�o�)��yj�דQ�i�j��ީP��H�f���t)��4��F������Z�ץ.���,��XD�"W���G��t��x󓸰�}�5���'��`����� @Gkgt��
�TX�и �DP{�ҍ��i܁�,
P�fI��C
� f'Bv�����:��~�sgH�g�֝����aҩ�N�s���~P�/�=�?���7���ϡ��O����h������Z�Z�睜�iq�<:E��3��+���'��<�p�fb�K�>��*��	Dٹ{������� �/殦+X3���Z��F��.pQ����{��YJL|���|��>��P��J�),}듡�X��M"	� ��V��S�Tme���A���P\: ��$z������Y���g�}.bs9���r-͠;�$�u�LXQ�C5U����֧F����l����&�x)2/��G���x����!�z&D��{�I,��-xi�`X�I%4|1�q椓���;P���f愤dPi��&+��[�����t����5m��&tG��2��!H41����LPT��
���Ƒ��1�~3��,4n��N�r��&���^��]@K�tTxԵ6]DԸA�貼�@���*S�CGr	|O��v4�Eo�%�B\�-�LK�C���� ��َ��ɞ����(	1�����������r=݂i��]��ߊJ�����;��V�6��צLO-3?���EF9v�[lkE����[n�D ����d.e�:��ܯ��'=ib����l��S�\��-5�x��{�=.5q����5;	�m���Ϛ�a������� �Ϸ�Č:P�6�(Z���*�yh ǿ�ń"
㷩�˱^��!���f�B-=o�p��BHY�i�|�?��^*g��J�mS	�H�讦���P�p�`	6Q�Y��󯞀	e��L�_D兝\���S��ǋ���H�2�R���;Yr>R�>����owaT�����l�1�P�y�n�2��R���O�wf�#r���p���=�Oj�����T�0C�>���U;T�q��"�Gl�)xd�>J;=,t�O���g�n.������u��V��?�ęP���"�}Cs�l]�4����P创(Ӷ���Ʉ�m��O���?�u��,$��2%ӑ��s_�����v�	�Zs;�m�ެ7����jc��T~��pD.O<!A9�"!M�{�����@Q���`������Re�$��w)N�W3�Ø9�M��T�ŏ�E�P�Ԇ�;�0���M�E;�P�9���8:��b&o�"NO�����?Uy����Bۄ�Kx�|@�:����2Cp�Ù�*��2B�i���ǵ�s3��D�	t/0[Ln�v�Q�ܱ������DI� w��(���hu<�s��Ns� \7VŽ�	���e�L
+�w&t �,?h/�M�a�y�MSA����{?SX��/����M��!��R��.h�F���X�H�4��t�N��_$вB9�).��8�O(䦁ֻ׹���E��AiA���썓�����Ղ�?8G���R{��� =J�M��l���t��Kz��TXxݾWR� \������}y��6����ݐ�f�j�O����ԃ��ya|Ƹ�0�pM�����
���8R+߰�:.� �x�zCG'�V�T�,���%�x�#=�� �{�Z � ��:���0[��؈�c`f[����Cv�+S�`Ё�hlD�~H�v�`�w�5q�ӄ�����k&5O���Jf�K�J��Y��,��eۚ��Z�޳�]��0���&�5������1;V�~7���ؤ��9���;��؈Z���o�f��y�|��o��]&7=��pV \�2��ja~y����2�I}�LG���L��iO���S ü�>n���yq�hmR��*q	a}I�vă��L��Ϙ�5WZ���5v��~������F�ʰ�͊O�Z�@��)]�3y5�h����t��\!#��Ni�ȱn¥�U��!�H��;{���{�E�*N����g���� 7�����\Y(��`+�6ϓA��ɕ��n��:�~Ì ~#��������'�ų]�C�:V=�����?�a;z�z�� +�B�(��d�d��yѽ0��/��F��6%��Η4?=�pd,E+O+�c=�j{�=��S�5 0�{��"��b�Y�ɰ%<
c���Xz�FL�L�W�h֚k�h�+�)aP8���E�������E�ۻi�ôtZq��y����,FuY����#��f@aQQ��n5��o�.�eR���S�B�:Q�h�{ڎsM�%c�� z��ֽ9*�U�[���o~�+�E�d7�o�u6�J7��nFIs��@zI�q@������9��x���k������6�$SDSjFa�����L}�,�L"X1��(1��Fo�:[u�U�ϒ�zf��#�6�~���C�9pĮ,=A��{�9�.R仱�k���d�O�OV¬��1�ln�r���@�;Φ�S�����I�u�[�1�뭆���l��kek���2�?K�y�|��YK�lP�y�n����n���/	�e莒���.� ��2�]7��a�k��:ϣ������u��Α ��?[�{T�[b��C�`sRt�m\��Ѷ�tp��hq�YXZ���g]W
q
����S^�c<�>�����p�M"��z셌1�M��v�w4�鴕I��MQTB7��a`(��_����y\�i��ذ�)x���$�D�|����:o
�*a��ݮ��=�T��*�v9',7���`���b��X���@,��ds�%9�u�$D�3�>TD�G�b��He�r���#�|�ѝYT[�k24�����1���:eU���C���PT��1ߐ8���%��t
��Z��Z���\���\�K�&j<-P�S�t�x���'����❽�� ��ĭU�"����ST�p`����+���_x����uF8i�뽎;F����՗{�7�{m�b9�);�wz����{2!Ԅ�-�4��m_��AU��Y1"Yi�.� Y΁0,1��id��?m�#˛�g�՛c��&�j�/�z�_Rn˶��a�Z�IwD�=\߇�H��o{�bH����
gC.E��}�zR�R���U �M�I�~M�y��{ޮ*`�a�3g�<1�_��t�~�� V"+�h���ȟ�"o�2��e9���i~gf��"��j]�)��
�d@^��Z�W���@�-��G����{:��%	hvg����2/r1x�%#���MQ�m�)�#0�w���(��(���&K�m��d��E��
-��q*g�p��0ύ1��e��t�H)I��R�[9�U��Į����E���j�c��X�Rc��ĩ*��R�Ϣ�C�Z�tqQ����V9S�$"��H�h���#+^�d7�@q1�����w���rE�o��ݠ.׽��a�a|��\v&����ɦR�k%E��G�)8(�Q�՞��si��2L2��)�|'T�D�J/O�]����L"��N/)����c��)�/D]��n�QN(t[��� %x\V��%���UMԫA˴���S�3�$��9�ľ,�LoG��m� �77.�C�w9��8���F�U�s��o�ǲ�w��x��ue���r��	+/�����y礻>�̨*�mc�F�=Z ��"ƙ�:!�42��!�����T�E��
��� ߘ�,,���a��M���W�Y�&H}O�b���=!�x$���ӂ��$j#��'�F�H����rR��fB�ŧ���@�t�`!��'��d��i�p��W����9̖D�l���ZRs��ɕ2��}H��8��yM��.���)c�q�"N��_x�
�V=%͗��xz9P�!L�+;4��#���<	�Dһ�j�%U4�� ^89�g��J�b L�ڄu�y<G�niׄ�n���Y�i��Y<���ݒ�k�;�[ �?�ͩxH�� 
�	t
��,����ɚ3QF�ݷuϕ����[d4�L���D�m~�3gO,�C�vL�w�f��9S�����	cQƸ��k5�����'rac���z�&�oLAw�I/pl����	���3_�c���j֌k��X]��1Ӆ�;�b#��e��aS#����<c�1�g^I���cz�^y��4P<ӝ�D�ʕ>�����"�D"N��/sL>��^+	5��}-M_��z��{������kE~��wוj.�"�B<�о�����7Aܭ,G���6�v�eťD�	\S5�Q�Z1+꺑\'s)���ٜ��kAb�9ɥ>�u��JX	0��-��qt�jl���H >�W�[#�b���7��5j���	���mD��o~�0h�g���b6"����l��6��w����"ݷ̓�<�d8/�p�[m��_��.��G@�e�����wG�QHS�:4�� �����Ӡ��念:ˑ��4j����]�y�A�a%�>��5��oWL��b� ����%E�pW�8啙/��6Q�W1F�$�jba^y�T����iWԋZ�8+Yf����*�
�9ڎ��&8!�b�1����a��1� �[*Kf�WKw��h� �����K�aU�4��%��9�v���J[��K���s2��c?�5����V��ww!�����"B'���)ő���Wgj1�>X��/ۃ
�|yl����#;���⸱余=�?hY��K~+���yx+r:@�9ݛ��K�S�Ȩa�{ER�)+թݒ^-k�#��x�L�s��L#X	�����M���QFG� I �-�c���m�}c!OTޓ͙:Sx��[�9�ā}�M��ﴨ|���;�5Ά"��""�|u{GFj���e�yI��T�k��̹wL ���>���P&��t(o�1�n�M���b\��ɷe���F�"�U�~�<sC"���\�e�M_�e���(���y���w֑�[�ң���љt�9���'o\��*�R��'�}�)�	N�J��OE�==�ݮg��V�XP�,�*�s_o�[j���ޏ
���MZ D�R��rX�ၛ�:�1�����do�9�Z�G�a=0����s�����|r��M|��٭��0�����Id��悦�H�ݓS�$T�d-V�ۿ��i��s��+����n����(g&�7�#�\E�x��4Ke�^������p�� (�͇V)�h��{����%M�s�[\QLD�a�T��-+���� A�m���������$��%&w	��]�B[�����c�qLл�Tkf�/M�dh|xQk;/�tZ�ީ^�z�d��=WԈ����	���ضIFp�P_�n,�4KN�K�[d����d�|Ƙ��Jo,V�h;�T�«�Z��?v�H�?�ْ�����7�� ;SN�y	��B�D>�AH=%�M�4�L������(�L�8H�>� \J���(�.��<@����� ��ץ�m��|��)�k�}��:�����r�&&��1�iQD>S�<����s.��cI5ǥ�0�f��d�/B��B�g�X�����W�X�=��|2W9���s�� ��Bt�\�5���lu$�s�2z��
�wJ�q��eA�7��҅�PO�4�m���꠆W��n�j����v��{$���wH�e�`QeX �al����p��ڨ�f46�j����������eyԓԶJ����oL���6��t@��	]��,�B�u�xo�k��:�<� ~�Cqm�3��L����!տ�~�����8�]u3��d�=���\ӣ=�i���\(V.9H��Q����i�{M��,"� &y�Q��K��B�l͎����i=h��gx�Isb���k>{�ܣ�<^�\F��V���h��5���B@��ʔo)���g;G��ܼ�G�sj*!Ch�^.ٺ�#���n>��"S��Hk8ޕK
�J�t�rz����h��.e*%~e��@�O�sl)r����I�����:��[J�.ɯ���=(�ހ=��	�yP7�uš ���0�i�k�u)Q��I�'H�Ͻ��H�K
�O"���?��0f���J@�
�*�V�0d��S
k��?V�A]u������d�n����
9��-�x�vl0�c}�9�}��޾Ч����*�N����"�I�Я!�c!�Z-l@s����)�j/u�U�xPeD�FA����\ģ���x�&�O�`#Gf�k#2֝���@��U���8�E?F�bM=[�A�� G&�,�3�[O��7-G�m���hì��:�`����m���f!?�`��'y�L$+��,�2kS��l��8��kvv-`Hb\U���bn���U�(�NZ⥡ ��d�k�4�Hڰ�}��IvõJ�u��:��[�*A���35�Is<����zf*ɹ$N[uN8�QP�%��/����t�Mj	�X��+˛�pi����rDV�>�`�[o���ٹWx����ĦI+�+]Glh��pQF��p�Iz����3�k�ݏ�[v.��jCu51Q�r0�6�����Н�x.	�i��J7U&�͝۳��	���k�:Nh�A��QςD�s�7� ���>f�=�Z�dppX�P��I������>�C�%���;�KD�es�/�VY8�H���&�����*)�X�8񂒼2l�S"�9@��''9���v�<n|�N�sy�e��r�W>�5��-�����7_ZŤ��䊀���y�n��^���%�"��zJ=�}�*�4I���@@�}~���'~񃝄�٪�9�И�s�V��_����s�iʸ4�'n��Xi�!ZB�� *�T�(	E+��r��^�� �w��vG�Gh�zY��5cp�����-ߓ��l����<|~�i;�^����Ȳ�K;��s�{�?s#t˳<4�ғyv[s<���v�w"�?��o�Z1gw���}�uK�^�nC2�i� W��	Q{c���`/�A�I���"��e����"�|��H���P��	V~vb���VH�Q'H���r��aN�������贁�ҩ�g�}:�7���&P34�0��Ȃ }S�@�Y�|P)��V�KX����ɸ>'E��wIt�n�)$(�0�V��1-������҉қ7.���$��3���ԫB$�`����g�9`����1=а5:Ip�f��{_x�UD��u��^��µV�,}�B�u62��C�+(��HX���8pZHݲvvd0Y"�$�����K�k,�h�,^��4I@�p�W���
{���%�w���7o]|��A�#�0L��k���j�� ��]�O��qDG���:������42D�i����Ƅo�ʤ��1h�<�oz��k���=��c�u��wO���z�T�Fμ~�![��)��3�8&iǚ����h�SWӖRʇ�ܘb.4�����T8��j�7���	M�f��mh�G`�>_��㘳K�˟��)Zn#!s�^#r.�g�w�\t)*|e0���lZ����X��Cq��b���ਓn$,�׻�A�(0=���m5�xmə�,9���o:JE�=O��9��ȓUՀ(w�ZO`��l��9i
/ALnʣ��!WĪ�U���Q�B>o�+���#̻k��n��5y��W'���LAڡmN��H�V�&���&��Zxd�':�>Ǉ�=�'u94�l�f9��@��`���H��Y��:�V�= d���r��y�����"%��r�K�3E���cq�U{���q��:߲�G�|t}��G@�_���4aeա��W���E��2�m�m���Ʒf4^���<�O��7N�O�c�ْa����n�����7�~�_&�$�x�Ev���Jg�Ov	���m�sa�$���r� ��@qP~Wp���ݾ���RL͟XU��o#����ii��jM��g�����h�3ڥ2׿j({�K\C�.��I5�@�f�9/�N+�f���M� o��S	u�c���S�����9�S�騖�4��jZ�M}�V������~�����շX���	�e��G�wny�{����[�@@�u��h�HD��
5�0m��ڣb8�#T���nX�ƻ?l[咨�^�Q�+E�����כ९IkKU���B�\��Y��g^��@g�(�p�m��SF&G�0 �����0;f��wY�p�!r�䯜����aj��3C�ق��腭��YKE� s��^N¯��{DQp	��Y7���K2Ʊr�/�8�7��f�=�J���|ps���&�Z��z�g4ij�?� �v�S�-�=��'Ib$Y�����iE+��l	x��"��~��gw|<
��䅄�#�F��z��,�X.��~���P�>:c�}��$�������v�p��U�}�j�&(~���zz/y5�V��*1�k5�_1\�/^7��@�G�}4*���<�r�P�����s~-+c�Hg}�k���?��l��`�>E9.�Q��%�(��C�|=vߪc�	����V����`=Wi����͗=��0�D���V�b?y����S���ѣXH9S�TX{��y[#����������:�:57��?�^9w��y���tV��n�%C^��(���0Nnj�$H�r��}[$րKs�GL/�3�P���ƀ���&���<4��aMt?$/g���䞪4t��Z,��6(͖_1)��rIS�u�^4ȸ��uXzM��v��{����k��޾�O�.2��&p]��a�}f,t5���H�d�U��Z�zh��@Ƨ�Y���/�T��(f�b1��&k�w�E��J�]�]93��~T�9i�V���F��[��	91�҃��˓�Ś��%Xݠ�Q*�S����$�"�nN�*}���[��B����(.M���J(B��X_I���xd�����)��Fv�D�M��T ܎Z����(���7��
W ���*B���@�:0/-W�?��̕|���qׁJ�Q� ܥ���YS~�բl�V��Hrye�-�4��	��* m���}����o�(:5�,-�w�|��-i(��E$�ִkQ�6���n�%��������#lS�u\��7�AO
i��;*�޶�o��xV.P7$\Ȱ25����ሞ�
�g�h)mH'����<�T{�h�t�_�W�d�;n��D�F���J���E����4�И�����Z�m@�XX�,��Ⱥڎ�DDnT�U�p7R�Y<A����JzԸ@������j�h
��S���tt���7�~��\�)�6��lz��h�:2��r{�cc1xM��1�p $��s4�lS�an�`�h�)�3�
PXA���2� ����5���ՀO�,yΉ�u�J�3տ����=�˗"8��"�C&�l��-�?B	�K��_DӜ�@;<�;�i��<�i�-Y?ʼb0���J��1ç�V�9��R"8yD�K�b�Dn,k��ŎIǢ��4f��y�;8��S�um{dh510�Aq2�m]���#����+0�1 �]2���K���LD'O,��e`��-f_��TU�T���.f���u�4��v�97��p("K,H�����y#S(��3�;G�W���>`��ϸ���� ��0=���<r��&cK���S.� ����V�Cs���*��AxJ�l��Q�g�M׵�#����O`��a�G���T5��d�\~�>"�m�v��=O!�R/}����HOΫ��E���i��:0D0�b+!T@��.I�tB�(��¡��u�V���	p�����]%9x8�e��x�8Ӫ�mxC�%�E��fs��KdCS��Xd�djr^c�8������*zUB$ܭs�����}�l�A��(�V�4dmnWE�[�W��Н�{��~X]�ͨ?���3��\p��f E��o5-�}�j��I#%����BY��N�j?�)x�MyG��J�H�y���{�@WO��*}%���3+�Ib������9ʣR���k>����@ i�I�K�8z����w#Z�|�!��?�<�Y�0g�%(ns/�̠�[^�z\��bqqtL�_@���/a�����Ǒ�;{���v��BG�2WG�\�t28�� �Y�ε#���1�gCЗC�Ȧ���8@ntNkf�.��B�;	F.6͔%ǭ��,Mw]5���o'�rd��%7��Px�Q���~"�c4g��B�&�)�%Oe!���.�\&X�uX���+1})Bnע���e�x>�IW�v��Ă��ÁqGemN�����M���pw�}q�I�F;���e��9|�/K�֔п7eL��uT�� 
��K�]P{�-~�<�=����"q�X�I[}�:"=��Af>Y{��P��AY��c��j�	�:!a-͑
��}�㮜�<B��t>G�t�00�,\m=\*���뜂M���������ko�#{� �O�E���4^������{`��Q1�V�~a�'���&��<V�/��^,�G�/b�E�}B5{q�O+~ �kм���;¤ZBM/�����b\�����폫�y�]���	�_��K!iQ��kߖg9�:���o֌E���@���Sb4��ᗽm5�D�PRZc��f^��c��(��r��̮���{�U����9r^E+�x����g�&���c�7��-C]Khv�uՅ���9�/3�p(��8^�_�-�Ұ/ɳK{H�mIu wh�!�ՁX��sox[�2�MÁ���ށ��rdC��j�X���ˡC����x�.���Gi?����8��hr�j�i/�.&��8b�l��$���o��G�;��Z�Z:�T�/�$ ��3�Bw@Ut�[I���0U��;���Ǔ6�_���Hf��keX�}�� n���S�	�$㨎"�a���N��Q_nPh��h�Ed���O�_��W�Bi��`g��F�W��懀��b^;�=���,1z�ԎU�'H�y�H���gdE�*�}���)d*_۱c���z]�$�
7RS���b�8�M����|X����L G�1i��,|�|I絣8A�7a�r>F��х���� ����X$�e��"j��瓻����d[N#�OR)�p�����L���g71v��¸�.�~�Gc��Ќ�-�4�	j�/xkW���� q/(m�`�C�:*���V�1 ����VNDQ��߹����	� Y����&ش��e&�a��?�'\̧��R�Q�?�a�'h1��j���dj˩���犅��"�و�Z���޷y��+{��kEI���+H$�9���j9��&> �V�v��"؁}�Q}�+NA��W��^Թ�~p�14�?ض?�tY��Cq��_WS�l�"�DJ�刼�Q!9��:��꯭��D�_M-qa���#���<��>��}�N���N�ͪ �/N�l-�kxY���_ZЦ��26R%���;�[�OYJ�k��oK�>��]�2@��!#�.�`�����]0XC�Z(�������n��7�;�۽0�yZ ��	,G�������I�}�{�QP&�&�:h�ӫE,�QQW�ϫi����U�G�XG.���#�,��h��m[���:�ӏRT�7]�z���\������v�1��,�/ ��G[#�fYѐV���3�|��cD��H�=��sг��Ό@�a�j���G�ط��Eh"3�E��ε6~ 	���������}xSfS2�^�3�Wiw��`?i��R����'k�X�����&��|%vc��<<K���g�+��RW����8��F��Ъ����5��	��E���CW9���ZW������v�p�6�	�r\��ė"��V���C1K���m$e�����)i�\�ۓύ>5��������U�>�uҤ�?��v�Awvְé^��  Ps��
6�,���ݻ �����{}=��~�<5z_�G@5���5�������?i��e)�nɤp<�ǒ��[����*���?�~��o(��ƒpL�~V��v%�M*s�t�;�ꥦT\���~7g�D	5/��?1n�F���� Z�*�����O�����$TJ^� ��n)�!yțOV<_(q��C��^�y�!��d�����(�
������X'P�=@��{�nK���˷c\���I  �_���&'���hY����!f>���R�n���@�H�4��3?�oJ�b@���9�<8.l[��Cv�N�.����dnSi ˘�x�kD�3�
 m���^ڽ�s�g�mqs�l_'Ѳ5���j��}�6���"��wK����]�N"
ދ����W�>6�f��AD��F���t���ʘ�.@x?b.�C�1�U��4D��ҵ{�Zbe���L��)�^��lt��m���DpQ�����+�jmL�+_o�B����~d[�ؖL���?��â����-��sM����=�7ʹ�:za�)������$b�\���g�d�}sI��czM2{��Lla�Ϝ 1��̹ �%6�ɵXJbwq�����*��8 ����^?Z�{`\/i�� �,B׉EQ���.v?�7�ǒ�D��B����~&���y�瑑�E}R�r�z�#�!����(��-�	����J�ABNfA�ovg1*��L���>�;�S�����$¡ʈ;�|5.�ďj/O��g]��Z4�9��P�M�+���%�gH�2k'M�+ #�<�����y�^G�W��C�襶ަS�-��C� c�4+'')�B��U�4�ʟ��(��o�E��k*���á��bj��fg���uv��;đ�$Jh������[l��*�ú��ێ��$�?p��z�q�엏����O����O�d�\�aX�Q�N%�&V��DT�/[�ͩbSzU��9G���6*��٣���h��<d��e�"i�iAbI�=)�a`Ә�F���+��l�/9��O�m���C�����a)^���7�U�@������f��Z0�7�}C�$�������9�A��k�]�A���`�4�mJG�8�6�r�	T�X�օ�`���]�j����H�1W��Aa[F�s����΄k�:9�Ym�hH�ǔ_Z%�d���3���&On�Pv��k��-�Q�.�� x�՞�~f�+�>��)�T`B,w�zAƖ�F&�Qc���`��ɂ���������kA�5�xf���qs~��?ׂ�3�6ϊ�(�(�>Tݰd�˟��������_��؀�(��)���y!�|Z�#�SD�fI�D�W��w�V��g�����z���䠺|�X�(����a9��I3�os��h5Q͚�f�k6��ǵB0ĆBa� ���45�if���j�G/�lF,�\��*�H�:{?���m�}������]���nre��q���.��ӳ�J߉�P���8��q ����fX�L�p5Gy5ѵ��7V�TL�� }��|�����"m�RF4:G
PP��8 9�ަ�ф�6)}0�*�ͺQ1���x��LS�'x��S��rU���jY��i�X�ߜ`��д3.�3s>�щF��X��`NT$�?�Đ�D�*���hrfŋt�Ioe֌�+3~���E}O~ȝ�������rU��o�U����D��0V�I�JatZ�>?��4���-e�!�oӖDmЙ��($#`����-�]$\�Z�-�n�Z%�H��U�����}' �?`ݜ6��J�Z��Ke�4<���ƪ_�1S�(N�X&��R�0���%��l?�	L�0� 3��M�Iv��o�:���2]��V��僋j��Z����	-���ڔ�>�T~�59�3����}yC��~��8��ï�%�A�^��k���鄩�b{�Q�[a����� 7�F�$(�|�~J1�6�f<t�|�l�����ԏ2�cF�@������F���DY�&	���Zc��X�"g�1�jk�t|m�'n5��k�k�.W^��^���� 4oP����tLi��J42W��d�u���G�R<-���J��ܙ1z<�Up��Ah4�� �ղ�A��9/[&��,H����~u���rIRغAh��Xz/����O�lB2C	��E �D�o,پ�q��\[����y�ь��H���D��}�G��H�<<d"ϑ���] eH-���{��?KKvqى�m��� oM���FF���;��jC�����>��A>�T����縱�H҃��>K�w��~r�>�b�V�]d���.$b��v>����l7�O���(���1r`e$h�(�{8�L=�O?��	��v�V������ �16p��F��D�=(��1~T9��q���gT�#�w��_�ޑG���ݾ�V�c�����>|��)X/6�O�NW|�l�4��_��p��C�y��%^�ŤuWo���ul�k�?l�Vo�?�"g��@�=��蚀cl��&r���8ň۞'T�p� �\м,��	r$f�ڱP��K�y�b�ÜcoV��ig���f���E5]j�*ko�u���ԏ�=���M�ѰC��6�$��?뙋�Yu6�ǡ�z.��ɖ���cSwr��`>��[��p���O"�Ӝ%�$�#^t�8Ҝ��8��SU`V��Z����Tٍ;*��W-C��� V-��W0�y{�Z�	i��F�~ީo�w�tR�W��GJ�e=�0��ϑqk^��n��N���Ǡ��&�z�#u�u>$u�E�ώQ����Q��<��~��v/�48�=�b'��	H�^�eڢ&�lR�d+�+_Qnl�!V�ӹI�ȡ�/:h�]l��WH?;�1�3JԗuD��������r���ȭ%Ma�F�h��^�
���Ah�a[d�6�\Cev�Y����P��1Km�ݙ%i�'JQD��u/~�O(�ߋv�zkM��4b��1p7���%2 I���bvp-�}�G��Z�#A��3g�h ;k͖_������Q��JLZa%� �{<�@��N�}D�m�l8<`}�ɫ��Lڤ5����@I�xK�bmQ�`���N�ϒ�,������m�.:c\����sRP��6L�*6i$�i��i����}�� �����[EH�iM�Ϻb��5b��^�������L(~eI��f��ἇ���C�Wtm~�����_�/�2����G�ΗjafF��m��	"����dh�6���A/�i1���t,�_�|�5"���fw���JPO��)���_
�4K���'D�.ŶBD��
��b�B��k�\5d��w2�Z�?(��M�Sa�P��SI��پE@Ş�����vȝ�0ovγ�|AIi��6�=+([<��?I��;��0�]}�K=�=��2�)�������_[ф�LO�*["oi�f��E�Ojw�=CGt���t�B3���+���Js�b,:��FoUh���ֈ��i��h����1Osm�p意D�����0�
+Cc���᪰�dw��$;�E&G��z��K��E�lw��C6�\������"���>���1���pw���ѿ6�r#�H[_�!��d�>&�Fo��č��}/�1�|E��Pb�/���4�a��l��Zigϔh}^z^�6&g�_����k�t@U<u��M��4�~�+]k���Q�=ux+�X����v��@���NY9k
���$��3�2��Q�@�H���N,��U�ԩL|�H�\Y7&�cW1y�O��H�|ݻ��?8�8�Rd�v���r<!f4�O�'rΞ7�O>7<�w�'/�s��f�/���.Ȣ�ԏ�W冰�ZU_�G��Q0P%"�jzݗJ����(��zH?,���9"���+��;�Mn��<�fY1O�����'h�� �Ӵ�2g� ;�w���e�;yEc]�{FQj+�xV��)��Â[r�BL�: H^c�Y���%,�k���{��hO����Ie�2��Ҋ��ӱ��JZ��R%k�e# 5h�֨; ����D����hF�Lrβ>.����(��)�$�(�{���[(�o�c�����vQ.�{��'o�3��Q�	u��bC1�@��^|F��	���a���Y����3��Ů���a~���B)�t��f�@�mW |?,�%'�nH���!����_�!�>I ����L���3���t@+dF�O0H0(��[�-}r�����L�9)��b�=7��/F��ȏ���A���`�%�uZ��/cU8l��p>����^
���Dm���Ng�
�r�G��HS&��)caò&RY�!D6<�U���i��:`5���@j �N���{1�`�p:0�-PCH���\�6�{|������������N#�Pn���-B>|�
U��)X��_Z?�AC�:����(�'_z��R���yڴy��� w�jD|���z7"�R+:����%ȅAz�O������wW�t��Q�`39���|J�pم�ա�\⑘]��b�3�\@�Q��L�|�u)�Ck��4�Z�諲!��<͏̟�!����]��AB׎#
�'����J���_h���I-B�,:S�9|��@���$���-������^�=�_�Αz�%�[��ۀ�|859���'� ��0"xcM$&��F5$)q���&��%��9x��Q��H.�(���u��ٞF���a�z/�l�1£� �%c���-��X���_��eD>���(���ͦP��5_)x�*Ӯ��V�B|���@n�R8H5�f#T��/#hyh�ܤ����@hVl�H	���6�_�f�a�
�w�xN.��w ��<U�2��A��r�'�I�CG��W���X,̪ʂRW�!���1���M��ݻX._�잩�]ؐ�}gSF/�84���c�x@E&trZ����"�����eږLL}
~��W�v����ƒ�E����5@I�e��X����ɂ�9���jp2`kY�qg���-�v���\jb	�V�)Q"Y�)��S�V���v�^cY?t��n���M��:������hu ��p3��y��
]믺4�"��;F�3���h>W�b�g�Z&$���֙6r*5=��������Sdmk�p�u�5U�-8�����oR�n��S>H��,�ƈ�޷~���_zE�-�ۨ�����{�Ť��l�{hw�ҷ�����Yv*���Y�g��{4ܗ�:�f���k,��XO��@�]� �y�.��p�(����Z����z��? ��x}��Y�	��8Lh�'���j��������v��� ��H�sN��G|�8�z��ɀ2)�a2ќ4@$3���s����Dkk�6o`�ز]�C�#H쀦�a�=xy��<)��要 �>�8�@���p�,��]��v�#+q/%��3>�ћ����TL\��kV.�r$+�g[1>đ!��W���wg���ؽ�I���Sی(����P ��}[z^��M�f�y�5T��۝Λ�R+%�.rh�y��v�ۑ;��
H~ɇ�!y�d[�p����k<�[jj\:�����Z��7�bV�bL=H���2� wӈi������K��$�}�n��,�|�0E�f��}��;m��WhѾ�8�u{���O�,4�4��2�?�a�=��c������\��"�b����Y�b�	Ժ,���2(u	H�pĒ�z������;X�ׁ!�B��q� ��)2:W��W����:f�I��p�Ma.�*��YBmL��l�+���x�Ot�lӵ��D��V�r���e�J��T�)d�*��e�Y��6�kV��p-19�\��b��{�CѮ7���t�/�4m]@b���V��
3��t.�@������̫龐e@ $
r2����}�\u|Al">�`wޔ�1�?�S�>�2�ɥ-�n!�	64�;!0�WA�'���,�����iF|�6�sņ\`�z�䥼x���e����rNj�I �k��mSslh�M��f�仨
N�� ٱ�5g�\��x,���(�>�� ��pY�7#2�|�r&P���i�Ұ�y��m^~���"�Q+�mL`�3�]RA���&�!��5�<�7��H"��j2��ЏC%B�Պ?�A^�k�յ���I��6��j�XJ��i���2�����XO�b�xơc���obB��޴3}��1�g�*F�2�km��`����חm��0	IZ~b���8�g�%�W���E�j�}��>"�� 9�0w�(�Cߞr�j�5Ա������N�X��I�+�.bOX߶	���_�HG|E��m������m]���6(�+h6���T6r/��<;"����[+��#�+&մ\�	���
#�-_W<!f�4��cl�ӂ��RFs2��j1wz�	ՐS�p�A�����ӆajVs8��X�!�gU��}������n�P1�e|��
�0�Z����|B�*g܊�db�B��*�TQ)·�fo�nx��e"�����T3�P����ƿ3��1>�ǄeKi�ҴN �~��)�Vᧉky=���G+�~�TŸ�{#S׾)��+��E��}`��eЈ�#l/���s7�R�:�J�6VjA�Y;��{�68Q�J'd�ݨ���|�D��n;�1���>J��ה�0eDse-i�i�*��r��������4�cf2����I����L��Z�澴;��	�q�d�s�LC�M>��D6	r���g��̽����~�U|��C�bK�g\�,?B�8���U�():S
�=����^k`�h�QI;~�9eo�u�CS^����3��y�~BW�v���՚�w
ӲU:�U޲5~���H6������
XS0��)����l�%�ZD6p�L�(2=]4?��Z)_�KY<zD���Ҽ5����?m��vܩ6���?"�7n�V����3�6��8W��A>�s�vS��x�r~���\EZ��:�9�LY��SVq>ޯ ���z�T>B��(ջ��6b��
��V��/�Cq��剻�V�����Ȧu�1�)1�x/�:�� ��is����H� ���ZZuCO��LI���|�xMLN띗��[��f~n�_к�v]�{��#/�#D�ژ�k�b�Ǎ��w�*.�w�����/���Gc�s��� ʟ�T忖��,G%�e�>�|Q�L��=v0k�S�\���]��Ժ��Yd ���o�X�sg����kg\�ua�-��>�Vǋ�>v�ج\�����]Omd>�'?�a��ʋ��v��)o�s�t����\6A�H�G�v��Rf�9�軐�V��
���yA+���S�n�K��=���uϾ�.=��XU�J��h6��y&Q-���{�� �����g^�c�6��7���<w��,h�jC|p|�݌�����p+����Z�����<e,�#U<�8
�ؘ�GN�{��S�/�D5� �J|�@Pl�8"�-����~�Ca��B��SqԸ�BF9ˤ�����d̺�b��y0��f �ܑ��mbQ*3���|���த0�[�Yqy/5�-!�0xB[�e��uo���dBP˰��H�xAy��#W,�. �ߢ�H@�j��~O��͊ly�0�����?�q����qp1��[r>�7�'�h;�d#�Z���d,o`|��&�2<m?/��-�hK<0?��Kwd�d���5�)���&n�o�'IΤ0 ��Õ�mE��3,]ObM_��K�d�����AM�P^&m�g�K�a��+�����c�uQ�}!��~5�On�nM�>9r9�MT0�ɘ����[�����LK��<`&���U��`�Q-Y˅�,���]!ɾ�K��\G�У�Im)�cթ	�/�T&}(PARM��^��	�G ��zS�ک$�r4��^��fgI���QX.�ī-�lNnަ�'��Xm��FՓ$����o,I�Iԏ�8 Ah�w�����dknW��k!s���\�;���t[/��a#��TW���I�SfW��8�섚-�K�_�t\/�{�7�%���ex���#���(٧T2 �Cm�1㩴��";�gu0�߇���8j�|�LP2.2d� 'w�z������=˗�����Ԙ��:��6�0^��X"�f�Kc�Se��I�k�T嵞`*��n��Vl�rp�x s��CUd��a$�8՞�|���_"+�#�����'ÿ�Q_'�/HW����v֊�a��������K�s�0���`aAVѳb�|�Eн��n�%@\�w<K�)z�xF§(�%�i@i��I�h�sss�g괾�˾��~(Ϯ�PN�j3P��ޮ��떠�V���!�l�̗���
:a� ��*��O�
A�q�^@�̑/����/��dA����(Š���,})J'ondC�E�7��)p6�-�+~Fq1��H5[!gOF{!�d���"V8�ER� �%+�snͧ����o~Ȕy��a%�\�����%�Xa�tZ�J�S�����,*���Sn��L�Ǉ~�7�h�瑹�)SƏi���ׂ�Y8]��F����ӯ}TJ�yG���8��,~n�>�x��K�U���qLUj���g�b+��wN�`#x�u5|T���R)!�P�ʴ��v�X����4��F�h\֙G��=���&6�E;r���X����p��Z�,6;�(޸���[������j�\o���[;V�W\��	'H˕��1j�y�=�vv>`iQi���!WA� h0�^P[[/d�&)���Z+?�d��y�\:��:st�C�ۤ�ci	t18�y���׎�{x+:��c�H��g�N|��g/�5�c(f���9���=N�]i�sUη�@�����<0pd�����i3O/?�S�:L�&ͥ������D�� s� �n$�t��a��m��� Q)ɴ� ���P�o����A�E�B;�n��>X�5�h-�/����H��*Q�W��>�N`�,Le�t�����H���8Ζw�I��E�Y�/�s��-9]�rۅ�z-�۸ر�4ڠ�#,_��P\�����Z�e
��#Kֽ��j4f2;���������9�1B�w��D}�9�m�Le �#���Z��o�M�ik���7�+��L����."2�ҡ�>��+̃���b����m������!� (Y�#Q -)�@�����6�0D	�1ɘ���&	���=�8�Ի#v�J9������>��~@�n����?,f�C��M�y#���%�&tF��u��NB���Q�8�Y�ݯ;����L���Ჷ6�nU6��3+����|6vU�كU�υ`��~��9(����R��#uwB���ZI�=+D##��s2O�½���?�g��l�qvJh�C��_����X������,'�hX���>��M��c��X������X��W�l\w�D�h��&�/�%��jvj>��+v�JH5�캧%�=�Gې"��_�-���ô��љ$\�Ar�W���G�x��w؋$/-|�ӷ=#����	 ����Ƕ����\	���?�%qdaR�VL�D��r�������w�\�%�%����k�l6	=bq*��R3����i��!�[�l������=�
�G�!<ף��i�f\+����L��e@I��B�\�(V��Z���%��ھiz�Β��B'5�"\�5VU���~(8��IR�َ��Z,�6"�<��}��a%���Y3[ T~#t���Cm6����Qz1)��ɗA�v-��e��]�'�'�w8�yүB�8�P"3��LD�� F	m�lq6�Յ��9`�Ҿ�xھ�{����n9
�����)�y�Q.���ꏓ%q�%�c����s����u�	��s��)Ħ�ӽe�yT�C��p�ל�����?8F��Y9�Hmb�"��@B�6#�!~��ž�i=�F�/}��fߩ��rV��.����h��ԟ��o�a �>e���aɑ�z!��<h�����x+�g�1�1C��sMOD����U��9��n���Fm��8ym�p���֞�G���\����x�Ir�d��+�6����c��<��m�p�,J��g�vK��-������ϥ)��\O�|0���%t�L|�IW�C.�4���2�'v�vZ˅^.��4���3�c�����i����o%(P^�#�y"�i�M#
AM-�[WpM���ʖ��%�.�O
1�����d
��?�'�Z��]����U�J܁�2��[��{[ ��j^ٰ��%��!�rg��!�1N���J��Yk�[.��d,E�˗k�n���y	������A��5��<�D�ؓ�ф�&A��yΪC�	�A�1&!��t#)��r���,c���8'�f����IE��5*`�j�j�DnV�m��_��������d6�!�q�g-#�Xs���`�k���ļ���.I��*p��Չ7�{��(r�K�!PVNSRڮ8���Y�37|�	>���G�yt9�Q�"�k!��%P��Ƅ|�_�5�Z�+�f`cE�4p1�O#m�`r����#k���Y�������	�3A@�C�rE���9��h�7qLCMY�'��@W�9�w5��C��Ѩ^�}��ޏ@S3c>�|W�M�9��zB�n2� `u5.z�n υy;�sN������-D�C$:&�5�
���'H��ڿ�r@)�"�xwR��hTB�M�J���d7?Y��<:��QN�X��C%����_၄�]&sʥA"S�ʆ��aN@�[��XJ�?T[���%w�,.��<�����wBF$�U�6T��yg7���~�0����gѵQ֢̣�k�P�h@p�����&��8��$S�'M����3(���e �Q@�N��q 5���(c-Tj~���sˢ�\��c�ZC��O]�J�)ݫ��E�s�0�Z���9`7]h��2�o�t�����/xK�����0qg�ϖ�񏲊�Ր9�m�`熽�����ھ(��p�����o~6�8�>��=U���\n�g�4��<��]��5Wˀ�MP���e�CC#�����X j�kbŕs�Y	O��ң�����1�v��%����u�c�����gSkS� T)��B�,>�O��$�hJ�=@/R�j"$ۋ�K��-��=����O��S����)v��g�)	ݵ�"���Ł�6:tt(0�c3ᯙ��c�C�Q`�_�`uz�	y��0Jmɂ8��)��x-U@v���Ǖ�-��Q�hjʻ��u��=>��;�Z�iG�o<�Oà��2��;���P�r"!�.�s?Ǥcy�P�b0��4����g��Y�b�Xu����X S�o�jb1����?AΩ诼�GǛ����ww�z�CyVΞe���Gj��֤hm_�ǵ;�Aޟ!�?��h4*��49m���E+�N-��$�t�������޻A/R[ɜW��Ρ� G��t��k�u6d���M6�_���n�J�p��'ڷ�ȳ0��^�A���J�m��$-e�J�� ,|�:�zZ@]����h��U�!��D�4�<j���ͅOvn���%^� "G�#�Chox��a��v����Z������2&�����b��H��T���6��tt�\�v4�C�����f{�$J�z���Csk��s��L$G֚��.O=,2La\s7a�/<��m�Y�����_U�?��ı!�/�|����ac|�C+�^V:Jm�O��t��Ӱ|�_�	ꔰ�p�0G�\��� ���s9���C�t��!ei�G[kЕ�ě���Qb1�]�M�W�+ZhE�N�R��h=��-�ӲЬ^Q>�.�n��y>�a
3r@^0�+�J�ԣ<�� �U�������ʬE��D�@XVNx�'�%Z0�E�e�ݵT�ܯ�U����%�{Y{�~�T
r�~��'����'G�����5�lѲ4�he�kaں�$d�!,��ֈ�v_~{D&3G��,N��
�_~8tQ�Id[�;;QA�Z�s���o��mN%���,����yBc��q(`�X���F9�:��r��(��e	39���f��jo�~�k|m8���I������UɝW�J����U=I�`c�jB?��Q�k���8����i4�J����-_B�H���L¦��/�����sS�+�nu���'���DK$�����	��RQ�e4r4ۚ��c^}�8<<�Ȏh�j����f�q>�B��y��E�/� �#
���s"u�2�a��N?��-��z�̌jH�o=5}��֗���+�-c0�d���A�����Q8���rC��6M-(�=����Wq$��Q�_��J�(r���"�P���+����Q�r��U���6M��atzOpI�������sa;�����Dd!2��Y]9A���h�>���g�-eQ<2����0$@��h��b��8 ;>y�D��r��>h}{.�[�:��삶�a��2���B��d�����d�ҏ@x��'��E�A>�F�E�n(�-�w�jD3�xC�d��M-���˦X�����t^G�V�)2|b���f�Ӽ���&/�c!�<�Ւ�@��� �X�MN���_Q� ϒ����<��w�SU+��JZ���s����.���J��X�5��-b
�����k�� ��ƒT�b����=
aI��� TtTM�M)��߻�I�s]�q�5�KK4������A�|��	��$��:7�_�a��|�>I�>A|I�`lϧ��qM*���.�I-�!��*�M�m��L8owmE��/`���#}�.|��#�_�v0�侲�n2̺d4D�Y�7����N��0�M�9^�!�P���5@��RΓțA����H5�������ؼWv.}�<�������(�}B&}����.�"�b�8�S�A�ތ��;�1Ϛ��^Z?���w����X�;#{����J���� �I!?�x2��#Py~�����D:�*���yIm��6/Ω�?n�ı�q��e�DA�ƫ�pt~�R}xj����� �����Z���o�
�-�����z�f� x������d~M�,�5�?�Cf�s'xY��X�f
e��0q�q��tbP�T#��A�C��f�����#�,�ºN]ڐ�4�%��C���`.-� �0.t��z�����9��V��|O-�l��S��F^J��6��,_�����}���t�G���"�Ͱ�q��[�$V�,z��U�O�+�R����V�L���f��?��F�~ �E��H�=O�m��eJ�����9z&q�`A��JȔxh.���;�������Sa���x�H��}i?����bM�Q�gy�@O��~)!L��%�95ܽk�Q?����3k�����D�_���?�v�>&(�P��^��SƷ$��*b�j�y���?�����T���T�Y5�MWjL�5~P�1��WL�&�NY���v7zD��<%�Л&�h�Q�i�%ǥ�C��hj=�@��Ӹ���U.M��2#5x�k�|�
.H��.HNt,�����_������o�0��;�``���� ��C�
��������i#�1s&�z���uE��^��d(|{��(�lz��,�'Ox3V�Sv�a�V�z�@R��T����0c�9��m�����5	���%�&pq�������i��="sq�B��vIt[�s)��*S��%p2�=��٬.�?p��l�^���	��7��t�r�WÙG�.?'�I{�:���� �r�9��|K[��ZG,�����KU����?�5�y��J��p%���J�E���ӻ!�2>T���Qشc�=� ����3|9��˧�ѭ^��JJ˻,�6r0��J����#���?d������q��ௐE���l])0�߹I�`��/C�߻�ډ��fF�1�p+яnTR�X���[�c�I�v�i��!��OL��#��ݨގ�d�֬ն!�f+�����f2���_�6dU�u��7.������R���P�ϊ�a!D?����H��8�s0�����81���mܤ������/�|�0�����
�R6�5)ԛ���_��y2q��]~g����xҋZ�XC�9(pbo�wI�O�;H[�n�C}\����[E��C1�L��W�W���������o�z���W�"�����r�j�3�B���0��D�Y�C�	Ė�<�}f��^� �|��!�MY�z��hUܼP��*�Ho�U�IK̓?� " o�Q	�o�j�h����Oh@��|�U�[r�+1��!�T��7�s%YF��d�8fu��KM�����	q�~�x�<���J�X�vsBLʛ���ʏ�J.$��~��I�i����[p/�m�� �6���w�cH� ����3E�c�#^/��z�F2�� �./(/ox������G{$��^�@�����N1����`���}��?���
U���7�˜��#D<qd�iYۈH�o޲.�5��ۤۂ��$b��Yj>"�k;���'휼�+:�	�6j�h *%��ᢽ���	ʕS#n(�/�r<JL�Sf9Q�B��`n+�J�1	��Gy��An�HTt�Sjm���-��5g��X_�J��K^���@V��m��_	k����3��]����9/���J�u��}@=��{��d�$��O3��@(Ź
d-Ф'1�[q3BC��V5K]>�ܩd�!b����Uyz�;i��� ռ���B��}`�,iH�P�b�̀���VP��Ol#��5���-آ��I��%	�ڗ����3�90�C!�%U	k�L;����t+�uI�FX�A?*<��t�LT��d4�BL���W�-"��W���Ԑ|�~��B4����w�u�W2)ʠ�r��nN�G�`���!fs���NG�d�ƅ_�3<y,��^���x��֦тbN\���U{2�ż�ɼ��X՘��jl铐�w��i���@��P4�Y��~W3�D���?��>��L��<��~2�*�%8�_]P�F�;��Gk�'F8C4�fZ��`��㉒M|wsR�Bޔ�_?��i��xc���ꗾ[ri��Ć˞���'՜�mm�/��<ލ-�@��r7�&�@$�r�S�l��cc��Ӿ�l%sB?BT$�?Q�:.8 �(�} ��z�7|O�ɛ�����N!ښ��y&�(�,���5�S���4�\�k�A�����,�@���qHQg����X�M�A���d�p4@��	fx�w��8�[1;�|_]c�օ���5Fk�$�{��8Qm��ʖ��g9�g��+�_"�0�O6E��J+��DA�&>�XJ����~�Y�G.Y��eCN�hϞ�n�0*I�X�����`�4B}D*��ϭ��'�E��44y}P�v�)we�G4_���;�Y�n",L)�K½�_J��Ɖ��ض��T�$�������9�_4CD��(��H!�W��Ie��zAQ*�)�����{��nSrڬ{����"��Sl�em�����M͊G�it}((b�����ڟd��)��x��F��	ށ*; )�3D���+��8�I���(����}�F��W��v[?J �bXG��y(Z���x��g��Xʭ[g����{��q^�6��x�s��^����g�_hA��(�c
���}����:�j��r��1�44�Jv�|�+̾p��V1��<(�_2�+�u�6�L��T
�J>��~�CG_��ν�y/�j�g J�.�#�{�4Ӈ\�L] �t42�j�=0�4`�Mi�1V��e����ڮ'��\��֍��'�)d��F�`��es�'��e4z���E'��V�]�s���Ur�W4����v<�ja�Z� Y2i	�]�{8�!r݁`'�*�3	��2��(=�ˋH��5��<�E��xe�	��vL�eL"��:��3�S�A]:�/5��:M�@g���J����m���%��{'�G����}�z�Hȟ�f~p)�f�Ș��ʐ���p��@K)K�ir����~9�%���G�U�j�����Ø�=�1������"�Uv�HH��Vv�@��s^r�����Fe����?{Z��xM�cg6^����fd�N�0�/WjD�#J�F5����͸�q�G��1�� ��O�5Y^č16�R���G��F֔�h\�:{T��d�� Wɡ����!�*�,�tO|\A���}8w�|�b\�e��~�J���X��]٠���b�r���K�e�f5r��k�[�Ȃ��LW�g#B\|.�S���c[΃_Ô��%��nS��Ypj-��08���'�#|SUz�o��l!�u�����C�W�9ƃQt�#�g߳��&^�� ��_;Z��:i��[?��:���$��{�j{{�-~[2����"��<�����?�2�`ؾ��D�­]�Fd�}������; mŧF��d�v��M-21�ګm�B4��G"�E��-��/��i�C���+������=���$w���j.ޚq�K~�35��w�v�����@69r8t�-�rbƧ5S�o%����Or;*�B��>aaA��
/0�V�9D�i2�/Jϥ�DV�j�'�-T*T��2�?B�-a+$�Fh�ā�i>(C�LDu���J����S{
&k_l��0�W_�1��ܹ'�ِ\Hy����t�6 5�)Y3�+������+����/=8̭V�p��,C����.��<�����,!���*�4��E�1�H\��Ľ�A���0EAՓ��=}\�,��-G��=�w���uF��e����8��3,���F_�Hv�CMM�ܽȆ/�S�[{WQ��\��6!ۍ�H^=�����|���M�P@���jL��|�κ��Q��#uh톫��=�WU��=�ME>31E��V�z��������{ӝB�[Q�JI+�gyc���C6��d,��Iv��g����:�g���J�
 ��]����%"v� �ޠh�aB[�t4XHL�hm�xk�����e���lk�q8�(���u#�6N(�J�#"}�f��u�`�c�{��ҋ���u3x^����&^�"6�5��]��������'� t�����-��AR&�s�\+>YS�HO��ջ�VL0+�5*��j��H��]?"9�.�g�L��j�®Ҽv��/W�F��X$m�e��/J��<Qb�|�,.z�� d�X��ə��y�8).��8]{c�Jxd�i�1d$Coo�\�%��3�?�D^�ڀi3��DrQi\�V�Մ��Q�$i�=��b���9�Z��JF��P�axmoD7.y��f�g�>D9���9��x9$��z������v��Sf�l��C��a~�者󃦯ɷ7��䫾�JA8�;��a6�����%�&�_��,�#�
�ks�6;X��#�rua
�80���7�a)�f��Q>5"T�X��.l��l�d~��s3k�O'V�������d�930�jjل;�.�޶����ϑ�;#��]�[�͆��(Z�0.�xi@�����I����!��Y�8i%֧:#t�
����=��MJ%��R�w&>��O|x�a��{R;�L�0��{�a�B���[o�+�'�~0��S.@�D��޳��� =�������F^O��Q_��k���]�h��<�O�q���I�qP��^T�	Qo �x��5,��v����e棸vI�}^H|�#��>�®C��������U@W��3R*���6M��$ 5- +�qSFbǓ��Ilt>�?��:�t�ȃl�:#`��R
��o�ab(5ȭ��o9:��j�ɓ�B�
fZ�W�de�ص���P
ؓ0>*ݣ�&����A��oc��G�{������AX��;�C�ŦX�k������ʬ=8��&t���<z�ͪ �K�w���i�<�O�MC�����P*�9�?��<Q�!<��ñ+����R8�xJ? �2nN�}�|O�mec|�����)JQK���X��G8m~o�iӿ�0d�P��h�$Ϟh����3uܝ �y�'�J�u�qW�b�,���Hd,���_��u#�m��Pl�4�	R�g돦t8�=� L��BH��b�ml&����f�,p~Y�ip��^^5Z@P�<�2���\"ib�O��|!��i�XkC#�siK�9c<V��Bs���k�i�-r1�ʊE~�$4͗�7��EYd��ͨ�}�?C�rL�{k�nQ�Š3:n0s��#�P����(+�.bu�lώߟ'J[�������l�w���x��m+��O�;�4$��
g?��`�1[n�����wt���x@ߨ�ڗ��=�YP��������)?#�%������Jv�oO��F�xw���0�9{�I�F�K������� ���ּ������hwsR�R{�5o.��j�cP�bM4e����i�"O�Ԟ�
\PFK�%p�V<�}H�~����${L�sf�w3�o��|�1�Ј��<Q�e�df?a�Y*�o$�$�'<>VV�􉝖ϼ)�^oJ�w�7�+�vd����ό�	���ؗK��G!�OI��\CD��9}�@���T\��|���W3��\�֢� Y���x�����pP@�k�a�p'l�|G��E�`0�BTX!�ܚa�%Yݵ���~Z�v+���F�h�~��4S���ή��T.�k���ĝϯ����hߺ��������4:N	�������A�^��s�"���B�z�H)e�����ik�]�:;zw;��?���"���?f��efoQ�GL��D�&}��ȯu����
ٷ�v.�d�a�����q�"�W���俋k|g�2{��Powr
QR��L��\V'z�O.�Z1`���$���]C� �	@�q��y�
�Z��vs�&FH�$���U�y���s\$���+��_ B1x���z s�D����f����w�ƙ=���J^��ag3��2u���*3�o�lo���;��2P${Qz�c����qnJ�l�/��	��`��䜓��+&�!<�.�<���|duh�� �����sFU(�b'���2�5����P��i��s'&���^kw���$�6ó5�۶kॗ��2g[�T#*��2���O��K��!\8O�Lt�=��3@fZ�YIN:�{���W��{�6G�B#�
��P.��^kى]Պ�,���h^ga�лod�V�^Ғ3r�nbl���NƹY����q��<��Ȭ:�vם��l����\�R��/�fY>�K~v�Y^�a^S��p��9o�S�#�m�J������X?gr;!+�Sh g 4�y���W܊������Ug���~�L`:N`�^�Y�G�Y;��_��ڷo��H]�?��7��[rR���.q�����?�0���nN��T��r��:}; �w�=n�����`�9�b���WEP�k�I���ԩ����v�-��3%���i�|b3"|���WX���j���zp)O�>�\UM�P���)&���?�Y�˩�$Gi��f&!�S�Qm9��h���;�j��������I㙉�X)tD�Eor��|���"\�+�f�#{��$�f���NwW�:�x!�ݢ���bQ�\�����7k��e�]�a����#���i85ۖ�,s���קw��E��CN�lz��|(T{8��	�lH�a�t�9*6�Y	�о9�r���Ӹ0\��Ȉq�$%�8[��6�o�'�Z���_�9�$�ɽ5�D�;���%_h[4�P-�.��$�q����W\�Rw��NA�~��
9K��YL��bLҫ�,v�L���fz��`����k=�j ,c���
�89u��t.s��o8��W/팄��_�d��'��}��(�2����n/�� �W�3�\CQ�%K��L�;�������ы��q6����1�l�D�h��������f'Z>��	��W���!��t��F0еٹ7³��d�����WP�x�5��x�GJMr|���ǐ�T�vc��tp�|顽�ݸ��!�A=�be!�E��f�{�d���1�7�%v�HJ�� ^�8~6���v�7��aߏi�`��Id���JٌiȌN�6��	�C0�i�Z0x���c�C=����h/�
R"�Ag�9MA�4s(M�'�&�Zg������8��������'�u�=�����;�@E.û��e:��	��� Zf˾=p�ڨOЎ�W	�cx��T]��vؕ�_	���E�L�X�(��ux���ǟH�s��$��(���}\NdqciE.dc<��^�����?n�|ryE�5�!�E ���c
v=�!��{P e�&��/�Sy&�R�4��e11�
�������G�kxfa�>���<��^�i��F8ӂ9��A.2�Kof�hgf}ݙ�78�B���U#�/S�{��!+ Ԁ+�`x�c����xk(��V�&&�%˽�m�>�U�!���l�.��?>_�~@��w�<�+���O�/lf4#�3�)g��L�d����08x�,!�e���5G$�� ���tv�	]s���je���Y$%�3[�f8����{��(�o���Eڎ���8t�ʛ��$ų����ۊ7�٢���D�q��
.�?4�~¯�¢i�%~P�Кk׮zB=�n��kwc�?O�&�K�g�%��EU�T��67%�gj"KXn����'{_e��l3�;G�b�ȿQ6t��Cڗ�ˮ��3��*��`�ӡ�a(h�&�H �m�.�Ga��˙��o�9�b�1Y�T�ݕb��ː�=4Wv��4�Q����{��3s&����5 �� �p��ߓ���j���mQ��{���"H�_4U����-�b I
N���+�d���+�o�Q��\���cuA�p��F��7cIN�vb\��'w�^�%p"�q4���4_<���ĔJ"�����+���h�Z�ٝ3Ť��8��_m��B5U��V��Q-��s.h+^,|J���4�?[W+�BsN��0��cpS�itݛ@�x ���_�S��r6-x�	��=~��8u�T�

%*N��.�k����1�lq����k�c�|t�Rż}�I�Z���6���_��,3s�������^�:�:�߶m������: z<"��k�`��U&�*�zj��9��jԒ�6���E��9�U��CG���[��b��d�vڭ���1�W &���G⍘��*7���A����#9\-������!����匓Z���aّ1
�.0� ���Iq��ļK�#������+(�~��.����<J�g�{�a=�����I�=}�#o��(b���$t����͡Z�Lσf_14��<̧hf�s�o��P�Fc�nz:�����5}]�AA���1��N�����j�ˡ���J���.�Ӏ�؏���1���M��$���9���:�޾��K�"!�VQ� ��=���TwaS��'���
V��qa=F��������$Xh� �*e�/�Aӏ�I���AX�{�Z�`�0�l�E���EPS��U�tiG9�*W1�%]�� -�r�q�ԉ���h�d�nNϺ���	&s�U�%@�j�#w�(h] ޯr'4x7��w�{�"\�:��������@�r�P���G'��C(����t��a{�BQ܏��ٛq&g�^`�����?�)����0�bV~���zBZ���Ns����y�X�v�<�ԥH���mS�f3���s�	h""�}�����ʳ����V����}�=���ͳ��m���W;����a �y]_~�Q�S%�As�׻d��W�<��'$�=��.��/�.�9W�u��j/bh�.p�.�aT5sZ��̈F�î;�kh��R�f��m�
���</lf'^?EB�2#��̵�����+��~x#95%�f^�H#Up���͊@M���q1@*����^+W��q>�X����qF f��	G	_�����6UŻ6�8O�В��[&���5+���,sR3���%���rY�MӳOg�����?ʍ����}���𷙣%U���% ?x�A�6ҤC�-�]ՙ�ģҽQ67�S������nP�ߒ��c��J�cbi�[�}Y��f�h鲶�*պiҙ7���'�{�9u�K�B+"�����Y�b�Y���4�	3p#>m%�F�"��$E�团��MJ*���0�~�����O�.6�˘̑ �Dkja�H��������I�'�>�tp�ݟ�eR��AhE����k���a��I��2̈1u&�a�k�	��@�.���#1U�@!mߦV��F7t��)�-2�͟#����F��*L��`:>����3�4�<9h����0o�o�D��I(~'_OIG�H�d;��8tI�8'pȾ�Խ��c��H>P]7Z�%�!�f���i��,G�w0�"HW�����Ts�^����16��8-`x8ccA�M>h:���T��1\/<f�kT}���e[?)F#/\)6ڷN���]��5��,��++�k���R,��@/q���_]�n(0M�i�md��1����GsL���"�u:y&T�@y�\��]�������ۈ��>A���Ky؁�ϥ1��C.�� ��wm��,�z�唛c^8f
�ڠ�6}]�	@Ak�~��_J��>\�t���iP�����X\���;�R�K���ȷ��痮�ʰ�J�������)
H��
�d���v��8l6��N�e�L��~q=�/,o "�G�qzI���w����T��<_�lQ����5���B�0���]����?<k��T��U�ҭ�%�+m$7Τ5i�p�`��DD�܎x��z&N0�L+F~*槣f _�Nlh�M�h�������!��~�EZ�gR����Ƽu����⎼7�n8��ϙ�!��-�L)����5�8�4�y�<p��}u�]xI�&Hs9�=B�Y��mF�ˏ��jr\��^��-�F���X�
�0� 1�`$-&k5�e5�,5o)wN&�$/�dB��~�0����۽�06���ߺ�73߀�����=�AY�d�	kJ0��36�3�*�:��X+��b����Y 0�[���@a>�=m�����U��Ta����
�C��a2Q�^Ϭ��pL�͟�1�m3.[aޘf���1�@}�r��l�3��Y��`!9���%�]��Ą�st�3-���Ogl_�?�4*;_�3c�f��6K Im
/��oX�_}�9�Q7e���,�`�7�,e�
enadmP��q����5�K�������lX�qh��"��:�eE RGFF�aʒ<�0�g�� �%є(H��l�h�!��k�ˤ�.8�(�@�R�� Kl��bYE�5%�G���R-pBW<W�Z���ݬ�EC$�Pq�^�ȳ�ka�N����r���(�,�b��`���֪��}'m"
f&���t��c�,�(򀒳��e�G�P�ʴqs�����urB��. ��S�6 b�EW�q>͐��wru��C�%���	Fw�m^��C��4��٭�z��M\	%T��Y'���^�+dP�8�:�A2����98B]��`xW��_z�q�MP�9�o�rt��+G��H�~�9	����>a;+[O
̝$����d\t�Y�j��O'�mr�.{�IU�=�ޡ2i��
�������A=�=�C�4��IvƲ1����=�/M\
Y���Ӵ�$���
C�F��+U���ssB��.��P�/�X����r���уT2ȫ��I�ӿ����μ��4":O�]���=�Z�xG�Ƥ���uN^�~��ۼ'�^\Z��0>c���cb�����~���]�Pc-j3��{!hm߻�~���?ߓg���gB��H��{ig"\Ŧ���K|�ߚNo=�e^�`>W�sG�� ��S��6u/���>q~Bf��@N�\�5P�
S�=EL�����zծY]�1.��90V�����N�!���e������(ݡ�4�\�ůXp<�*3o�_�IPmά�^C5z~%b�`����bC��DJ��?�!(�*JU1ǎ�hS(N���=�WBT̕���]��N�g3���Ћ)����@C����(HI�t&�t��1�t"���IJ����(H���]]�췅�$2ח��ߚ�ؕ��N'QuZ�2L��K"���Y΁k�YB!�Y�^p2b6�l��W�~�m, ��4�y��m`������i$�R�+�f�/D)m"���}�UY���͆N���&�[�7��@�˺���sB�	����%yؔZ[��e��>�|��Yɠ�Aҏ}����\<��l���X��
�1H^����2?	��HN �������%P���w�wz"��1��즡�O�H_�~�Cn��5���s�����ߪ����D�f�T��l��=�&���CW��:����xF�A6"S��}��3X�G��kd�t�	տM�L��pڠBP:��Wi�]abnH���D���P�I"�`��Pb�
h�C�I�9b�h�Z2%��~�S8���$9�,�
f f0�B��:�6k.M�b��;�.o���нſ2�����)��č`�6�)Zt��ƙkh��F�<�1|")���Q�����}����a�G�l��@�,�97��P����_��\R
�S	tڂ�bd���K�V.���]�1Ե/-!�T��ŵ �p$ ��M�_�n����
����	D����U_�9�σ�=���9�PvjS�(�����
��oA�*��Aۗlu5uV�7���hh�����JF�) 8.���v������Z����)8�b��c��6P���䝒f����ҷ��91�6�>��.�����]Y.����"�?�8���;>KÈ[�Q�z�b��N\5Mzq)�e�Z
���9�0.O[�41b}L�D��?��W
/T�H8Bm�\$;�����3�	��?�67�H��z���I�:͆	�U�I�z������'2�&$��x�ȴteToYXi��^�6��a �4�Aڷ�tJ�C(x�ב�E�-���D��BNj�/�/��������p7�TP���G����lc���F\�B��
�ܒ�o�T3�a�]u�e}�-[�ae���%�+
�������d@}��\�s����΂����&�2)�����[(���F_�� ,t�f��Au�=s�%/Wם�K�t�M-��ބ	�Im��qQ�mJk!,� �q��C ���7�@dDeS��P�����W�	v�	Ɨ�x���F���F�!L������im.�F20b"������ַ��cf-��6���cuAkL��䣶�+���񘰞q��(�p�C��]�� 9:���Ѓ`��M6�����}�*h6j<�4���<�D}�#Ƣ�8;M�41 [/d�fze�4ُ�ؐs�_���:��׀~��L:/��:|K�*�\���Ӏ�2�qR�!��� 6;|K�[�SԸ��ih�	�p�FԌ�p��PȢ��mOE /���b�T�7T�����U�W��߭��#`��<���ű ��=���[�(a���_^g�o�KQs6Fۦ�Gl;�Ye���uȚ�a�V�bHg{K,+�����z;nգ+>�W��)>��qY��K���2�Í�]^|����Ѐݶ�y�U���:�UnM�4|��<s��z�(� rxz\���q�;/ka�w�T��&DI�\��|ϥA0���`ΩK�D�"A���^q�@�#̝G�6-����p������~se��-.b�����|~^���T;���2������m����k1��Ec*��l�D��8.(���e��Cq�~���W�!^
���z>����J��	H �L,�TZ�,v��J�j���nS���s%h;��H�ղvT�8N����z��q,1y<],2��'��@���0d& VN�N�Hj�<�V�������=�j�O���5LժBU��ݱ�!�1ws)!17���o�qqlg.E*�dI���B�T#��3�3rPc�uX7��#P�u���m��.�@���o�2���ĝ�����y0^րt/76����yj�٤cz<<P#>�O[y�e��FPZ�?���8��t���o����+��N����K��m7 ���}Q%C��.VL)o��T#��!�� ��o�۰�����SWd^BR������&�f�b�����Ŋ�a{oԣ�0E��ʻ��0m�.,�U]zM^�������@�})M�A�<;|��6�'H�5(L���T������C�U�H�C�A"�k�zgJݭu��4Ivh��uY�%�ĮX��ت�I�Y��}5��,`�%t^]A썲æ�DZ�K3���#�C�z�O�a� �>!�����pa��Bm/k��n�� eIS�ɷ�Jנ<?!�9���Vj��\�T���!O�%Y(�i���q�E�YF��p�r��	����j���]8 ��s���а�0�Er̙�����E�*ܘJ��b.ܵ�s�o���s�e�:�G��jȠ�ӣe�}-�m��b�A�m���4>��P�~�@�{�+V��$T6�A)���h��u��Q=�a���Y�vt=k��(�E�����+

���5���ই�d�J�9��X
���ځ����Z���J���ٰ�W�	�����3Lp�= U)�Qm��>�$����*��"�*9��N��8�>�\����u��jz2�A�1�,r�RZ{M����C�ħ��_����{H��d~�N���;����h����I.���ܣꣴ�(���4`��J���;$ǟ�q�Êqﬣ�o]�fѷ���������:
ڿ�T��_����.�n܀U�͂�Q�:A���w�8*
ri����ky}.�#�ei���N�5����hK������@���hR3m��ӻ�K���ߐR��A�`�|=Z���� �%8��;� �`'ՇU[�z����VO���W���G�����s�G�f�S߳�d��\�֭/��n�s�VE�j�F%�^����m�"����o�U�r��{�~���T�,������?H�4�Mz�6"�A�|��%�x<l*skd�����O"�������;P��B����]H�<�x�[�#ϙ�+��	�]=�hO� 58X�mpO����	WIS�}A��s;��� ��6�RRT���L�/�3<�;9E�k:��_���ھpE�pQ��R�f2��Q��͊��)�1���1J ��U}�M����]��v���>^�+d
Fq��Y�S(#��3���ڈ,/s퍃ďM�K�,w�_KY/��.8+�	�"|>�$KO��0�����5���4���b��F���QI�b�H(�RK'ͬ��Aw)������϶UH�T��o,����A�H�	�(�e��/�o�.o�_R��η3;FW{�D�q������b!_�|'���(g��R���Tj��ю_���~��^��m�r���,~�p/S�<��E?�e��@B^���/���~����1�?����V���-����׷ϵ@����u� y'�e
*x��^�XDWQ�Ҝ# O�qɃS�qד���v	ť#���d/���Ώ	�y�V�=��J��8�H��$��c��)�a�ރP:Ѓ5�(ڝ����N��N[W�x�����.$;�#�&T
��q��7��3�J@����j���79���fl�X>��KHL�֐߶?�ED�}��Jf�
U��մ(v�$���g;��d�ϩ�\��}֋����=��BnRly/Q7Jn���pqO��lh��q�n�Hщ�?m3�6.H|� �h�^R��`s2X�A�g_�â���>����D���94o�.�F�|��މ�SƇ�����e��(��_z�Ս�sYkl 4��>A�����[[��@.'�J�������E�gv�F<e��p����
�����������շ��dk��3��JE$vbQ�Tt\WRS[��Pg����T8��-��3!��,o�?R\�?*��K7d*q�o�����A��-�}8�߂z�	&�"��1��d�#$�.H8t�:mb�%�n��]�|���B��M"�u;���.w/N�Y���'��ql5f(y�t7��6S����gAtYkt�[/b����ڬ���_�}{P0���[��e&�n��m5���ȬE6���O��������H�0���K0�k�.��3�Rw�z�r��a�Z!=�q���E�q�f��}'ч�d>��R�Rq�+��5��Q ��he��h�]�y��B����<H	I;n}��p����ْ��"=��k鎼�؄�n6�Rp��_<��^�3`L���e	|Z}�QC�o"��a�͢� ,I����O�R��L�*��o����V��ru&�+ÄB��b{ݱ�)/��� ��M�OB6�K���K�"�g�xI��u�r�9�PY�FpW{ݦ�N�Z��/�Ա�O�f8Q�<���hl%�(�#�)�؆5-���^,/77-M�bӠ�Z_���X]���5��%#��;�PL�>�������ڗxI�|n� ���؈)�?Nn�B�WU�7kZ��Ț'l��c�7�q}I(�k��J�t�����z?Q&�S]d����֢��c�l�Js�<$�����W��H�AЋ��9[���	���R����w�_�9F��jo yl�2-��r#@ޕ/��͌������G��A�I���Dk�P5��[Z+r�A�CҒ���S�~�}5���J5����|�Y��y��������Ҝ�嵡�Լ��'��w�$2�<��D=��x���w�2+�,{6�j��3�hnhM0�W�"��O��s�HGq���2�b�C�X[:U.$;f��L�o�}�+���C�>sjP �X�r�y�o:��h�h��#,�̈��}�������"�Yw_���[�p��z����3�	�:.b�߅k�?�!���g��ćE�{��	䕭�FKD�Z._��l,1ed[լh5������hӢ<d�N��DӉ]������<�<�ƻ�U\�JݏY�֩�=��S�-�ڿ	��)kYD�Ih�3��!�,E�pu�O����A�`AT�/΂�D���)�7�|O߹Ƣ��4+=���)��:��{�!��#�,C?��9���H�q�bz��e�LLtJ���h6)��C�_�3l�a�����e�=]x!�1�>#�F� Iޡ��:������g(���g���m�_�� �O|�쨀7��U���ųkd5^�WSd�pou�h�.(-fh�������蕎w&nu��}��PZ�4 	��A-�<����Q��=瀴�d�u��g�O�ѧ+�u�w_���i�㭠�_QgU\(3���94\����!v�ΖP��V)V Ej�%��'u�E`8Q	�x����,�&�hD1��0�h���>�g�i,bMJ�b�@rFC���� ~�I�^c��(��}�ίgQ�B�p]M�l��/6�h�S�����`�|���Z���`��0��K����;��1��� ������do�߅��ܜS�h���זO{hlB��3M�څ��o��G��d������[d,2x�����:ӏv1=��zҰ&��_��<�*��N�R^��)�����]C�uvE��[�E������oE��[���)������.E�o�&=:W�{�L��f��	"O.)�uq�2�j]k9���vZs�%��ngvy�ʹ#`	��%�P��su���d�6��f���c<�^�"l#Y��"���z)��x��t+��O �P�uA�;a���B�ާ�ˁ���i��z4�F�"2x��VR�L��^��� I��Ef!��I%�0�{���g:r�;�ѹx�����`pk��@�� �r�4���N��ڪb�WQh|��"�<=̉&vۏ�B��Q����S'��k�����6_�C��PQ�R�Typ��^.�%-�X}'��됂	�Pj�;�a�Ft%�l���7M���ge]bx��:�BY|K#(�;c�'(w0I���=Ǣ�BPR]�]	��s!X�0��N-U]��TAB�J���,Y|%.�يn&�RAB#�����%�\�-�ٮ[�!���N����z�fz����arPy')[�	���l�&TJr���R�Qq��/1�ws�k5JD��ϵ͇:��N���茲�Ao�G���g�`�t�"�tP�����@-[#������Z( zL�o�FF�d�/^!+�3ԑ���!�Ҡ3����R�6�������d3����k��kM�e��b<%_��wE���ޥ�
�31�����,����3\����"Z��>R��u��iDW���ʶ��U�&�@k�w� ���������� m��Q�~ŉW���6���Ol�*������ �L�0��'#չ(�c-@��T<�Ksh_�x�󅹡G��~]I�Q��q�X	��߻*�#Z���@��'\:}ɷ�6���`5e}�p��d�@������]����ٸ�-i��"^�I�Ei�,$~�i?���ƳЪ�EN��x,i�h�az"
����PH��,{����g�8%+#~��Y,_1�z{��(��QU�Y��pա�T������YumB�4�o����-{��y*�(��2s��A_o�5���v�ߍ��A�H��h���Cm���B0a�`վ�i�.�YUS������T*'A�L�s[aoqK��T�:V1HP�ƽ�q�z"X�'yWN�Lw�U��Nx�.M���1͊H܋��w�C��s?��_�Ԙ�B6�f�m��/
��H(��i`���v�o������G8jWbWl�a�c�u`�{{\�u����']��=�Ո�C-��z�rLd�_T�X��؋������]����\&Y�����> �89cQ��L!(�j;vb����."�t��rb�F�u,G6������4��j��Wj��\0%�m����5X4~����o���l���W�)L}'�o�0-&���0\"Qb8;?/_ ��;���CF��C	ɩfw>-l*�PP	�jI�qe8�����QS`��"�~6� 	�-o����~��r��_r�y��4$@ѣ���~P�6�΍m/�`ϬO_��x����*�+:�-��b��)�����n�c�鍶�i���K�	�+�����ΡsR�#��}&c ^��mfpE!��|��,�N�0�!�N9�dQ�	��d~-���MZ����c4?B�a~��r�搥�j��OB	�aq�	b �_�Tɝ�0c:y�TJ�J�X�heĸ���M�v��7�.�)/��:D��-��1y��[#M��:��s����(���j=+X��ʕn��_�y.Z��ٗ�j���? ��G^X#�3���+��N�Eer��n�sI:Ԥz=�D� �ԋ�Ƴ�V�vo�|�m;R�Ƿ�ށ�1�?}���]��nz�&�=�Z��H��/�w�BP &md�.�	��"m�k-��D
����C�]�6���Ϣ>���e�nO�>�#X����q1���4��5���7�\  +��P��Ho���U��HC�����g�rI���}g�f�0l��&uIˏ�XLigj��(<��%AHp�,������C�"��$z��+	�@:}�� ܲS9���E;�_��}�C?$I���Z\�w,ͯK��c%K���oG�A΃�4@#�4)X�A���C{S,%�W����ʹ��)"{�����F�?�f"CM���-ŻsW`|��D�*��ټ���v�*���Y�Qg����h��ܵ�3�g-e��u-�Ϙn9b�#oz'Y�tJ������J�m#X7o�k��Ŷ�(O�v�^V|;4��1���-AWm2e�5%�A����eC��/�K�jb2��`�9D�������j)Ҳ�R�0q����4P��w_|eR]S�CV�͔e�f�қ<�-+��*��C' �1�{��Սm�I
;T�Æn|J+5����D�L��Sf����M�k�U��6�4�(��t��v&������0U�:�ۘE�����x�26�Yōd�I���rkP�y�	�2Ǵ�d1X�<ښ��ǇP�@�D�)
8��7�~3,@�Xe+~�!:�_�mO��w�i0�4�������Z%�8�Q1�	�$�?b|PI��������,,y��@(6�>�&��N�����3���~Հ9�A|?�p	���!�r�����1Q��}�U@Ҥ͜G9�����N���i9ӷe��M+�~�o�m0���an<2k��V�%}3B�B*n�ֻ�����ZIkD� '�I��{�l�F���A��D����yj҉��/�C/~��|R'Tw~��W�XC���þ��EI��������EhQ�s"/��۹>1�;9+& h)�C�����"B�G8M����=���J���m�|�:;����A����C"��`n�JS�h=؇��9�p�~�b�B�{vW�������;ۧO|��~���TB�\�j4K-X��hJ���v���/(7�ծ�ZP޾.��*-�5T�3 �_�j�:��2�bnxPNw�j�E���!,&6��1����0a�-�i(VB�k��"�Ϋ�?%�f�����d�����@ՑNb��K���IE�`�����\�OX�
!���럈(爋��#�7��:��H�׈m�\0��ђĐm3X�䇱*��)rkin�|LRcg�}�T���e'�����W<�B�O�ق�N/;%=i|���'������	�}]D�t���e`��zR��oO��yL��sL�́��,��5�B'�nB�����~B�3MF�|��R*�@Ea�C���$of����V4�y���Mw/]Ǟ��_|I�qB���y��5;��{/������ ~�ݻ���rH�6l�C�K$��5�H��)��_6S���t ��wkk��DG,�o�h�h�n�zl��/��YMĤ{�H���>�)Z���,�o��.(�α{�yT�?�F;zң_WB��;&<��ou�'�'Kl���pR�8c�.��9qv�����~����δ\`�\L�eװ������{��c��ǈ|�ed���?>����kq��#x����͡u��f�ue�oǥN؉���u>f��fr�$�8#@ #�ϑ$W<��`�E����N&��B�Wx\4���l�]7bHG�^��3F�q�kVV'g#��^n�����5M����#��md�釆m*G
�w���qJ{�>/��l��b<�=��`��){���,����?�]C)�P���@|/͆����l�yb��u����؉��L�)[1�,��9�tkҡ�ޯNwix������a�J����r>�*�d����4�����^FAUJo�C\�e����%:X�|C�G4Hs\`�񹌶����DeFE,6x�w�� ߒ,�Ɉ`	ߏi�.���V��)�l�z_�4N�N�ij(�O������XßA)���gt3TG�WK8�o~���'��$ǡ��Z�3�ě�I�������7������~{܏��z[�7�==���-8bȄ�S�톦ӱ����%w�呑��c��G��We2dN<�����G�J��ݨ��'��'	&J(����}�L��N�Cq_ⓡ����0����>�i<w��~o��ҹ���!�fn���Q�9��������>w����¸q�>�Ik�ƥ2�0��&t_�3���/1��4S���]����#`-�!������<�Kٛ���`��״�����,��
�� �LY�o$+�Ɯ}WX��zh���!��}�#��ӴE`��dq�N������s��	��<ȸIo:�`��G��Շ5�� ����������$+���\im��5����i�
��zS��P'�i�^@��*�n�U"�w��;=u��+<��3������^����aЙ�  ���B�|;D}#4n���$u��mP���mE���X!	���Y'Ndt�&�rY˟J���Ƭ���Uɓ�]�<�ؐ�m��sd�#\!)8�-�7ʧ�k��ɼ0A��m�E�{a�U�9���º�»yI��Y�b�7a�5	����V���B��Z�%��$�Ū
#:��*݄������ETƸu�z�PWwYp�.p)����7j�8��O�T$���<��\����>܈!�K�*���k�>��V�Ѓ~�I��ǻ�x�Xg�ϊA�&Z؃�`v�_zM[�5/Ӯl�U�z{@�b�����g�O�2��06+sR��?�ma6(��Y��W?+[Lά�/Ɠ�6�_�T���p�zS�¥t* �yeA6��(Dk �V�X�Ruhה�Q�C�>�`���/�#�k�����C#�G�Ϋò�(l׻4Vt{s1���X/�WQ� WT�<U��n���۞-������į��r�*X�����E����Pj�j�e�����2��<���o���m'�F��?	��0(���⬾[�ʙ�5o�b8�-���2��T@�G�R[vs
�8��9�ÒW.��N�F���C�~���L��48��C�й �1�Aql�xUr뵔�>L�KҦb��F"���Fΰ��*�qk��jf�y����8�ܕ�k^�g�����B_«�<E< 1i��
��Ν�'ym�� �������
���Ifv�_Ȫ'�&��r�P�N��	i�K0T�P���l][�R����0\��/��~}S`��xv��[��-V��Ȑ�L��>�6�v3@w�2�C�>��<֓|-�1��Δ5N�>�#7��H=l2��/�#X"��{"d��{��>��n�&�͆��mT>�d�c-��4*���|̟��cA�! ��΅z���>���@,��@y����0ak�/��Y�b����QJ+�W����&Z`.�<�����,�ʄjF�v��#`��v#�@�Z�Q3F���
~P��x�Dđ[����a����g!��祫�MU���^W}����k!�(�N�T+��.,����H��S1W��)Cj����{��������N���sS�<E��Bi�~��
�C}.�B�Ȍ$�7��
n�Q��^��|C~���.�|&�SN�����Bٖ��3�V����j�(���5F1RW�-��4j���'\�������E���g�#�	4�D�SטmpѶ����ݭT�(�2 �ߠ�$��yMuP���Gȕ{���>D��AV�Mn�+�,'�!�la�,��*x�?IP�Xe���ԊO3�Gd�XԸ׶�=e�囍�cY���W]���-b{�)mqs�M���9X���	��)B^��Ⱦi�Ǖ^Ed� RS��ۯ�i�f X3�[e� �f�<rt���A��ٕ̜�W><�Oo$��f�V��Wxs�^��K�)c�3��WbE���v,�3p5Lv܈�&�ܥ� �m.H$����ŕP	j��Yｇ�/RR��^aN�E5 L�<�5BU������:Grӱ�g�){����YY$�ԫHyI�|�Oa�ޙg�l����#2٬�<�,�s�	�?I�T>h�a��X�����5|)F� (j��uZd���po�Sb9����}�Ɨ���ͅ�w��6���D�b�us�Z]0e��Ql����q��]���+�ɘ`ȋ�8�Y��#Qr5�ɔ�1����'�������P�Z�`#�˕�{��&��"
O|.�o��^�,�> ��=���7k���!\䗐����f#���BU��0#J���t(�t��x`Ej��a�Q�S�?��ڍ���b\"���T���۝�i�%������m������B)��;>�?��[�q�G��hEw]�{�QW����Pὔ�elT��Ǡ͐W.>-��8��I+t��f#T�4�pL�s��nX�K-V��E��܇�pm����hNo���R�	v�%�D�T?ě�e|}((��o
��{+�0n0�����Z��-�[��ț�*�{��*L��-�|Y8���$_�f���K�<0!+�}p,2���"������0i���4nz�Mk��l6�Q����.�o�+z�:���������No"U�uO��U��ֿ-\=m�p ��"J.eﭞ�H�4�˙�-��u�8�k�h�`jה��,�ƺ@AB�b����������3�/��d�W'���hM00��n��uE���g9|�?PW�h*���Ȳ�9�ڡ?��QvkhasQ��!i�ѷ�H�����]�F'��F��OE���%��f�n;�� GR~���$w�����m<8 �Zvq.��g�Qԟ;���Hv:�E��m�qyܡ����B1��+�N��|�CC��_.�Z�-V����ǂ����j� 	\�o�E�ۨ�;����@ط}��R��k9ΐ%]3��]�Qy�����$���Q;Lv*@5a%���ll�^��2ߥWth�'��� K�c����eM�<�5nh_���"1Oo�_Zܢ#��PYl[7^����)�)`�H��3t*��#���#5��%�TPkrJ�5�K�{|���ٵ�e4��0=�*P$�Cp=�>6����Ë́E����અ��wwZ�6���&T�����-��n�W��a a��Y�2ʠ'�Y�K�f�n~XD�U���6Yh�0�j�$z�l�:�bl�e��M��)��Lݠr�m���:��;��ʕwP0r�gWD��ӳ4$�]��YW��A~�׆��,�	��=m#I�-_�8Չ��J����VV���(�#����=����O�Fΐ����H�Th<��X�������r.�w��2i}·�4��x�1a������q���|!�Etb�c���-0�N����'��^}G��*�t]�4q\_=00SVު�Ѫ�Qn+P�=�(�� ׄ���?��<{�U���t�c�$_�M�@ ��#o��R=�_�J&���g�p�|5�@1��Ҩ����� Frnق=����϶��Y���r�0(h�Lf���� `�r��n�XJ`�Φ`��PO�� #�B��{z���.������|��p�?zubኰM@_��olģ`7�d�t��5M�Ͱ5Yi:��1��2��\/\Y�g�!W��a����d��h�\���$�p߮������ �=��Ͻwii��i�`Z(RH��������w�3I� 7)�T�ᰇ�!%Z���<�`!O ��d�6yj�yC����؝��݅7�L���N:F,�<�Ee]{���q�'���"GunV^���FY��HqR�G��!F����}q���Y4�;v���H�G�����F�JK�Z/�<LV��U�2���dgt����̚PtBn���M������LL�Ž���02�����"��?]m�A ����	Anν�XC�	�z��8ݪZ]��[�@&8���*��Ř��$�#�/��I���F;��e%e4õ.�X�0#N���~����0|(E���/8!�</ �j��9��}?׊-"��f�wv���{�!C�Ř�t�8�?2B%!@mW���?Ȳq	�1�D�Y/q)x.u�����[b��9�.��W�;�e��|��2��)�-�R�2���:����
,�!*V�+���L<�}�mA�O�	�>7~�i�ts�t�4�k=�����]�|�[��� ��2�&ήc��6������-Ϗs$=��#��&<ߝhd��1c��N��y�x���m<-y�8�!�	.�i^ӆ�8(�v]#�|;�򵦢c�\�7ר,$=Z F�e�0|R5K��������y2m�},��>ӵu�r�ٛ�5�"=��%��X!�mt,K�*�nTy=+�+6vv�|�lt��L�!���,�@�~,,�f>AQق'�$>O$k�g��Xkh��c2�:o�ݲ������<ǜp���g��d�ժ:P�>C��y ��X�J�Cnq�_��
\DA|���X9���o�T��3hU"�&ݽ�+S�6[9�mƊ=�C�E��8"� �ȏYD���7���OT��S:*�%��Gd���#�CSs�K�m$���p�;V�]w��^�x6!�2��$�e���K�}'��%��L�:���z����.�����@���j�C�����JJɒ횡qd������\ۡ��K_ؼ+5�a=��;u��>�Ka]�͍5��D.o�)���ty�U� �P�Jm�ϐ~���Dk�ꑦ�!%k�o��.>��d�X�YZ����|�n���,�zS;�p��xC/nCR�a��Í|:���A�5�495g����i3A�V%�?�g��{r���������ā,s��%���&,c�т�&~l�;j�����uy'�^�}��s���q��:�ݍ��U�7��T1ts(��ӑ��#��J��]#������uT�.�Q`<�ѱ cU������>*l=��x�����ҳ!%`��M�y��A��Ț�&��	�5�������	��!x`;�G�c�h{�l鶾���«�-��p���!�M�O)5=�y�,�`b�x�{[
[c�n
�L8y��08����$@�8/���J;9�*i�����Sl�g&Ob��.���4U<��A�/�6����V�1�zP��t ���g��6��F�}q��(�����G�Ƽ!��D.:����Y��Ma�H�rXX�"���y���
�l|J�׎�Ȟ�Y�6ex媋�D.��GE��?��\(�+I �/�ˎekk|J9"4��y��n���L�4�^^�������X�� ���Yly �bӔ�����a����;�gK��g�0��M���kj�m����)��+��J�X:VD�(�T�(�Uʆ<�>�� M�4@ep�ci�+�N�/K_o��S�Пv4���Kz�	8�ٷW�jI�[��Y��A�̐ԯ�0����� E�5L�yDL��7}}0xaK���y#r����T��LѠH�����ށ�/��dz�^��ێ@�K�����49�K��8%�8����Q��;>ǀ^[�$0�e���HF��`������.���Q������"��˭�Ke1�ɓ;TۃU~����8���i�::8��Oʞ9T:�����;�/�~�%u`Ë�JgL ��J���;�
[ئ�$P�Q�s�k�wRYT���VX �~�>95����f;,6�>�ɿO��s���lɮ	S��}�ģ�͋&��5��%\��̀H{)?��]J7]
����5;��|7�P��[�P�:!�\G��<��yt��>2/)G�O辐!�E)���~�T�uB�[��xY�j��!H��F"���Dv�|X�d*O�.���U$$�4 =�6�'�?��ѣm|�>���4*��B�$1�@�=Ё�D���^Ѭ%��7!��e���c��O"�#�b�1t���%������ž�����W0�@�΍ԓǹ�不F���)���29�w��S�A����}D�&)r52����w�a;���&9�U��<��°sh��
_�� +����$'��,Y��!�^^o{8�U<�T�fX#�	�B���3��iyC3Wˡ�EA�$?��3U������A���pJ��Y��}ہMJ�7auh�xygf .��X)+c�;v.'������u:
�iI_^��A?�ǝ X�+���.����|U�������^-�*̙Y�����u� �$�ʻ����B>����45�Ȋ�
-Y�A�������4c�&��3o�.�l��1�� ���u{��mu����/0ń�Xb�l�I\9�����!;ǃ��Z�✉I%$�Q"���s�4�6޼��|L��:��;�y�m�g��w�a�����phH��"�>bQ��㪔�q�
6K'#���K?̍&ν��gI�M�<���+�?H��F���sG��2d���ُ��	�[{4��%Q�%d�!���ڛ��B��F��AM�|8�,��\�F�#�Y*w���	�lv9:��?N:�W�y��r:�>��3O� �"`�������E�������T<m��"��f��m�� r]hd6tyF�A�H�	1�͇.�a�qy6�;�D����o���h��g�X�!ϨdE췘��b�ĭ�<�s ��R״�Ǎ\��S���q�D�
u���?�#̐|�H�e�F��p��E�a��'�[9��s;T#[����|�����[��X�G�`*1�}P�9�79w�޷'���{���B�O���|ې�p?�7�z2�Ķ�"\*l�+N�]_��@���2���f
��v�3H��O�Y��I=G}��#	�y��k��U�H���f�T��xQ�m�	����:��`M��XT��Kk�m����`1h��Lg�Su�>���hM֛���Vf�Sq7R�z��8%ɘ*`�橏��cG�y�������>�AS=SU<���~��<9�C��>�UNeэ���E:K?]kM'��%��r2L2 p��RL�n�� �v����ߝ��{ؘ�_5/T��=,���	�t[>e�
�Î�X�	�zV������Ŗ��<P�('�	k_�=��!��
T�d�,H�����	�#"����M�lP/Bnmzq��Ʋ����c��D^��ur�H���M�Ps�촺�����Jg	��M��`%D�߾Շ���2?�=�]%�7�ID�:�!�8��9��K��4!4������ݚ"~�v��^��Z�q�[5UY�d�&{���,*ats���$u���4S�S�GB��˒���͌�^&�K��9�T�-'�T}�$�WU��+����z\a
�.���^<��>��?ʢ$Yk�VL�C*���+��ȅ�:��50y[��٨��.A3L���B�X��EW�d����?Z�/���$�;a��<�|5W�����.%�������U�n��Slwd��Y���xQ��5FW��=���+����Jr��n��%Ѩ�ŝ���9D�%8H�� 3ozEk�C.v��m�הu�X"�a�`�ycQa�_��|{��L�a�Nܩ��]�߶*�8�0U&>���*�}u�qT�J�����|�P����(���h�jI�tƺ핉�6��-p�hÂ��F�b���V�P�Ne�����(�hu@��}�dH����}i�-��[�n����w�q�n�#���.���z\F��Ě�K9��~�0"'"��f���ĶA�Ԯ�?�(�\����Z�͖'�n
ɯ�TE��R�E?PsLFbR�_�@�@ܐ��M�*RY,�A.��&�� ��k(,�YG>1��I�:d�
��<��d���?�����6֮�����x))��i��?ON��n����7�!�h���g𭠨�Fˏ�1�	s���X�|(��m���[�	i�<��,'k{wN!�E�|D!��Ԧ�I��ː�R� *ƴ����~S�m��_i��/���[����P(_�iVۅ���m"e�������@-ZƧA��š0?/���Η�؋��)����Ȗ�$銦�f(��d��k��/V���v��5���N"[,�I�T�jA��I����5���%GG,�:�o`*�맛�	�3� �:��	3B_��ZU�1r�B����qv���$+���:l����wo���.� �{C "o�h=H�x0�F� �p�Db��.}���Ac�L���+�v�^h�q�y@7�9� ԣeKD���k�T{HaK�pvu�a���6�D���Ἂ����pO�Υ##�qO�o>�`�>J3�R�I�3��u?Q���M��	xe%׃�ȍoxrRk1ڱ4��x!����¬�1��QΒcT�Â�?�^)GP�U�q�ʭؠ���3�ĕV{6=��r��,��y6ҁ�Z�;J��D3�+��^����ɡ��T�MN�l�}`�Jy����Xp �Q='������R�c	��8�Y�q�����Ǉ|�ߝ���4�릣8�����D^�5��8p���':<y��w�x-�14�kDT��.�%��Os�B6�LܰV"$oSN�&8��G�`�w~�f6��������;bo��:t���ܦ-!�0|i)����S~|�i~�"�W��î�,zƩn�B�R����u����a'��d�[��"#l��v�����s�Z=�gQ��0+gۢ˓��~K݁�d�KD+�6t�C�/�ac���`3�e9��&F�	\,țE|c.�U��'��սQ���Z��F�� �\Xpj�D)t�
�w&�fW�W��
��w��kBg�q�k��N8q;�_y�I�2-��o#�t�ܷ��
n@\�S��H�4(G5aMO4��'(%��f�	���{�B=�ɡY,	�$�︗/�(���n]^){�n(>��y%�D����F���$�l���),-��s�J�q��.�Iy�@y���0�M�B⁳K�US�À����â;CȮK�O���X8�� ��V��s��8/%̨)o�I�IݛY4xGf��>���|��������U�!��K������H��N ��nX��z^�ybo���u�D��S+��Fרn	��)���ݤ"S*��Q�Z�x����Bq�)���o��Ͻ�{�/}��T�7o��9���:D�(��)�{�T�_��a;�6��z��cL#D����9nb�����/��Vj�a�7#�Q竀���/�R@�M�
Ivw�6=&�G�K����Pq[	�M���@d׮���J��Y|��ČϜ�~Қ�Y������I�V� ,$_��2f[�.?�4'|%Z���!Nb���q��fSc���y�N/8�-���;�d��eڄ�T\k`��p�ǯ�9��Խ%��u��8rE�ۘ�8=�$����C���JC��a�*�3�Guy���oRj,Ҍ�(���9�F�Kq�MY^�S[��?d�$b-O��z9h�mD����c�������ڶ�����E�/�
�e�SB��=6�G�B<Ԥ\��O�n��N��f��c�'�3�@�z�E�3ZL�b�����*�.>�!|���ӲdV..�	IbQ;p��b���#~a�'�Y���=ƧP�&�8�E�a�B-�Ҏ�M&�R�:�1r�RË�!��_�r -���ak�1)���
T��TO�U��5x< ��ɢO��
�^���e�<u'�M�ݟn�*��5F�y����/�g%:m�A>��о����t��yڜj'@���I�F��k�����H� �n){�8h!6Ͻ��R�r��w�
=����4�i][|��q�;Pk5��+G�D t�����$���:���@��r�+
%;��`A�Iص�%����<5 ��.������5{n��Ӊ��qΫ���m���ƪBO�r���K�}
����,�w�w����H��7��r��&e{�����'��xO*��++�Y��	��O���6:�+cnyt�,^&x:�e�UZ�q��"^�z@%�S6U�i̔�ս@Q]?�/*�V��ZLjtw6B���HYuL��m����[ʬ�ۨTS{\V~��h������8�8�c�DW���i�]��Gh�2Q��sM�MEj'�!'}Հo��Q��U�̝�#H;�cā�;'���k[0k���8')��t=E�/�o/���w��_��ĵ3P��L2֗3��2&R���a��.=�5<
���K�f�bwd�q��P��� ��E�^M{S2.� ܾ���<R��`�i9%��t��P}'�5G����"��.g��ǘ�M�8�(��M�V�-%t�;�/Q��b`�	W�P6J4�6�O&��;�[�Ui���l�<C�H�yY�G�ED�|!Q����^��]p���ہ��w��m��X"_R��(M� ���s��b}K�4���2�=���K��6�L��B��Ѯ46� ����ͻ_��;i�E�`�l�Y�f�t���3�\���y�`=O14v�W@U9�;Xɛm,s�}���l.v��q_C+<��lJB�`�A�-���ÆUt����Ni�Ӫ+�Y=���Z*��h��ư�be0Z��{��@�aޑ��1�F�7lXsNXP¦d̄��D{O�<V�ܧ�_��g��OM߬=*৞���z�H�}^K���A8S��}X����_�d�u2�(n��
I5��vrˇ{�~Z3�HRi���m��E��*4[%!�S�;D)�߱|��y�:�5��=>���!�J�4.�,��}f�O\>�%�%�68�
DP�lLi3J)��B3Y��Z:�A��#8@JbcOrw�h�_��z^�hd��?B��VI�^���$�Z�%mڑD����D�>�Oa5m����m��K���mJ"��E�/��0���2h��,�`������p��B鸰M��ވ��K�j5n��d0��?E���ԡ��ԡ=L$�����>+�Y�LA�O�0w;�ii�wm2�ḕ�]I?	f���3������r}j��gduR�CK���߼pq�k���t�]���Z��
��4a\2V��"�{5��C�Z�^J7���������T��d��`���2�9�˿E!l{3��k����9���	��/]�e�\5l ��4++Z8�n pU�ǝ��Ve9T՜�-ɺf Wt����ʻ����^�C@�>[�ȌQq�:�[���5�CB���0�7�7@j*��{8�ul�{mwn��n`�;�s��/�O����EK=�W��j}��c�Q��w�����#��;�	��Lv�P���H��L��?�������lq�/�^���������������g}󾭏"��ܐ'ޓ�}V�ze��޾lE�X�����9��y%B4���_�%�mp�=J��TO^��.-�oz*G�?{t�Mƺ�H��Ys�)f���ßP��<����iLg�8�vin�N�ʄL�f2R*"���i�n��������y�S]Eu�ˠ�˦ǘ��Z��PC�$o��GK/zZ4�N���֬�r��c�7v}�:��XL�'F|`�a:��}�\���)��׭��nQ�a&E�Ņ�#�^K���4<�nO�����MM��a�<τQD�Wf�zr��j�|�	`GC���2�R�����'[�E&�����p�=���26>�7ݘF���d@�{�����&e���6m3.���L#�6&SΆi���%�[���K�����n�5�K�*+438ҫ
�sTZo{H�����S���y���7K ��_���w������ ��U�ݤ���W�瑼!���>%�e0CE�$�d���G(�����@�D�����%C����Y�vJJC(����?����M�]w^��s\lM��-���ݳ�;!��Q_O�����Z=�qpQWr�����̏�ėb7+��W�`�%����ڸ���,C�}��<�J�0��V�ٔ@�j������,%��"@���%-��f���ѷL#�<�񏣮lW8���S�2��h�h�:RUȁ��N]�	�iD�;���NX~'�``�Y���!�@�h!�NI`(p��ړ.3X�cSM6U$�h��~�w�fL�O��S�z\��1BQO��x|{i	�7g+-<Ҩ����r��cf~�7$�o(q��u�V"Y�n�P��Gʂ�V����4k<�@dG���P��5W@i=3���:�4Y���EI+Bj k6�n�pSy)s;�}9%N�[�B�#n�?a*W}���H%<((�* ��s�4�
Po��h�kk&��zu�?���u&��'�ֶ��� %("q��^����P�dX���̚� ���ø2�4Ú��clde���k���d@abP��l�e/X���drM����n*=�T/z]tM�����Z,�u8��k�`�-��s:0Z�Ïe0���7�QNE�4{�)u������X��X�؈��:ݡ�h���Է� R���c!
��~Y�a�Va��k��qxK����Ǫr�g��$��>��Ds�FO:^�������+{z{��۔z��W|��6?1��<��l&�#+����_v2������)kT	��������F�e�|z����5�a}0�a�.0���k���'�P��R��wt�k�p�E�Ć8t+�ܼa��F����jvC@zE|Z��zS��@xg6�,���d�Gm�u0f�z%���24�|,�Ҭ���	k
�k�[�N8�kU+UɃ]B�<��%U����C���X#@KΩ]A�T��+��"u#s�/dMS�1�vw��3�r�,_b �h��v��v"G�rJ���t,Q�E���;��ʙ���#L���|B*��VN1��L�;�nܕ�/���4���I���A�e��
4����>ծd����g�DPn���K�va��~#hv���k-m��=���`�� V)�����j�;ݥX�	��JI��[����ġt�u�/R��T�}�[�kO�.F�F��m ��gw����d�ҩ���h9����:��U���>(}������j�G���xY�n_����1eAd��B�T�l��5����fdМ�OU�n�'5�Y�@rQ��:Cֈg$���c�������Φ��5o��B��
 �ힴ�^�"̍Eǂ 쫵�@�ʜ1���D�f��o�I�u���xL��*��m�K#��%'x�?'����./�y��3�Q��ب�HV
�yZ,_J��A��pw ����f���t�ln���-������s���et�\p!�1�_���C!G�H,=2�\�e�}x���z58ǫ�����r2qZK�<�����Q3��.��8�t�2��iĪZg�<�C.���kD��u�p��}��/I����l���G4�����Vȍx�Z��C�,L��C�7Pg࿭"����mC^�'R�=z��Gv?�P�����ߟ��R���hj3�sV�3��	I�d�U��M�7�x<����ǰ�E����F��A��
Y-���hNie�� �iO�e���Nb�GB��k�i�GAe|t�V����e,��sp����"�>h
gQAOh��ڝM	ٺ�9(c@ٜ/0ժ����V��&�#��ɧ5|�U��?�0昡��+��rt���u�u���fp��P�}Q����މ0�t�@y�Bg��T_˖��}���^���2���G,��ڃ滟q��C�9���������_[viԱ�:Hn������pE���HJ��r�i�%Ρo��?-@x����t c^q%���`��.O���I�A�_��"y>S_<Q�ӹY�j66
z\fa�����%i�z9Y|p�	�d=}�;�Sn��M~l������͎*�o�ځ�{�@��<����l���.���K����2�$:�J�$��s��PU*z��+-`���o�4�%9���h�^����<��ƺ�
�=��v븰�y��pg�\�$dbc��=kFX��q�a��E�%Y,
�[�Z}�1�����2��Xt^�CヷD��h��;X���C�eC��W#'%��p|Ɍp�Ź����g����	X�F�B��hy��պFۖK�x`�y��
ȶ�Y����I��j~���� GOi#�l�*�Y���9'�3ClCR��<�	jhy�>���Y�m���E��}��7|�7�4��6<1�p�P ��'��:-�t]�C����ê�͠��Q��n@0��i
0!6��+�G݁y��F`��d����3?���c �J���KK�{B��ٿkO9v^��M�ە�azF>��;%�HS6�<�Çw,�0.e3V �h9��;�?0(��>_II(�H��x�T\ɼz�8���Z��k�C&�ڢ�C_|;�v��r6.H�q�?8mɆ�5a�J��'f�d�'poܣS��,����X��"���fre���~-���b����������w�P��Lz�Nܖ�ܿE��j��M�ё��]�~A��Z�kl��sB�?�Z����q�G�#��GOf����
U,c�%c	�g�}�^�OG��ѺZ���M1��~)$�*�(h/FG;ͳ����ؾGq:��G�>����Ehޮۏ6a1a#�YkJ��!���V�v��7�;�g`G?f�h{�k�ء� (n!��Y���٭$59��Wd�ٌ���<˅mG�ϋ�<�2;R�|{j9��~�!�#�&rt�xb�F(�v��U��Ârt}��6�o���t��`����(y���JΛ��0��KX��N����w*(���&�ֶ�N����z0"}��+2؃�r�gsw~�>-�E����H�Jy;��YIU���;�D?���9�;p��������%�$�6��%��ӑ��D��.�_.�UK?���G���ӄ[{Eg�YxС�b�Ő���A9���0[M\e���_��E���]r3�:k)����8��{�D5jk�1� Ë�h,,�~�Q��:�(�0ej�P�g)�5Q W�ϼa�.���J�<jn���)Da\Ȗ���� ���H��eR������ZC�����J���(�7Ə]����y���_��Sy�g�q���N ˁ���nu?�d'��9X�.���͞����\o�����):��-!hq����{����({���N)�����~%����*�� j\��&X�ᦠ��8�/��M�Şv��{ɰ�k�)mp�^m�j���*�>�l��/e�n��DuK9ol��?�w�N�fH�A�lx5?�ꥐ P��%��o鱩I)j樲�ǯ؟ON4�V����n��%�����؏I��k�ڊ��N	z����6q������I?�L�(54>5:h�������I����k��Ŗ+��2zN�[�������)u�x��>Sfu|��*�,�����5�`*���(bL����%��2?P?����˜� ~k�~a�Nv�X�;��J�Em��`N,-O~U�è/m�aF@���]�3+g�qv�&���9s���ӟ!����Ð���R6ƴ�/B��И
���7eW:�̕s<jݷﺋ��gs����#�=�u?�
�Sbh�1��j�1��XO�m�D���h�#9ec�L�qY=����	�8��Dn=HƔh옛ϲ�(��?����t���J�>�x������N��͝/|J��xD&]be3��HE�p1�WM%p����'<�Zt$�Q�nɆje�.�fr2�^��6���"���v���9��3҅��������-���?�Wp��$��R��4w�)O���ԛ�{W۠�UTDh'��.�è+��4��U�>�$/�YlW@��z���L���3͛�cT�1���ְ>�P��@�6� NcfS[-"P�S��;��k@����0���%�LM�7��)���gP��Y�ӧ�M����v��8�]\5�R�p8�X���5�VXQ|���T�6��1����燹>�oJ�U�Ƣƣ��O��C|����G`׽�Ҁ[������D=��T�3b]o�<�)�۸l��R��kD�x�l�XD�I˯��%w�f4l�,)|3����>�g@˞��*舟h�d::P�㶄0�N����w)�70��N7wK@D�F��$����X֬8�#i!��Wn�'�:uE�*(å�����"_�29P��&MG���4��:��Ȥ�u�g�5�͎���E��Em�jS���*��_�`!p����8Yp^������/�K�jW4aa��ٱ*sv�E[���/�9�]&ߞ�h^`�y6��d&�X����B���W���c�W5������LR0������Nme� ��KW(E�G� �Z���!��pO�,��������d�L���hS1��:�j�>y���(��AW�N���09������n���x-�
B���ܠB����Y'!����=�דM�suh�z\��evcbiN�����F7$n>�v�+��K�33է���d5 ���f�;scl���ng���7CoJ�j��d�*�p#ҫv5��_`��I7+�G2滢�?qDo�$H8p�!_B�3��&�50�_#8�;n�V��P��g���j���a�D8������$����AW��rS~u���+�.KǨ�8�'n�}4���bg�|�[���-UT�٬���q*�WD�bQ��h�����	��$�JΛ@����S��e&��yZx_Hh�х:������؁��	@Z��=�}��u2\�m��S0�`j����b]�$�� ��d�bv+�&�x�|N畔��)>_O��@���5��>������y��S�f�9Ӕ�"v5�Z�G�W��L|k8A>�WL����A�����c�:��+֪�-Rd�c,L*V�r�����Zo��x��v{�)e��7_��`��t�V2��&�`{`����^D�F
6�'~WE�Z���^a8�;���'���
/=����>!qg*�~t�6�p��������w���~?�R$�$({��J__���ŻK�x��!����wO�tPu-L�o	-c��"H�3�:��ȟ�e��U���T���w��!sٙ��D�T%_�V�6�l�."�@\~�YB1w$ʦ�G/*&t�8���}�w{B���i�z�[��5��bLg)V33|9ӣ�Cy���"����!�xn<���a9��Vh*������uO:�e�rI��{ap�r??���Q�*Te,,7�S�]���y�Մ ���vU�^�rN��{�:_�:�gT��!��ڥ�,�&��uyJ8�픭,��Ed�pN0V��$�	����׽��êԆ�H:
F]_�o���n_���^��[�b�B7�:B�r�}�Q���.�@L	y�έ'U9��;f^4#�}�n��(~���L�`C^�āb������Bp1����aϮ�A��WLnҜ���t�U+���~�D
9��ס~j��%����J� T��JD�w���b�+K�����1?�R����q)���	���9B�t�9D_';e����n8s�R.���f�jbL3!���D���s9E.W�J"�������̿yD`�ڌ1()#w��\� j�n�B�A��Ӷ�����2�Ⱦd� �_�%� ~���_��Y����h��8x�s���뒍�4[�Λ��WZ�Ji,����Y�	f54՝6���ۉ��������~'�����x��}A�y�[JX+�MLlW�.g���,1G%nYn��zvT�����0��?
�����?*���^�-JPT�O��������Q����V@�'X�]��0���b���cg7�.#"�>#���f�'�L ��(&K�ߕ6yů&Z������.q�D��ɏZ�$���읞� ��;FH�Iˍ߂���;�Y��{���]:Dhg���GJ�y���>.�Kb���1Ζ����X#V/�oQ�;���4�Xr�O ���۠g~$6�5d]�����M��*��/�PG�@8@?5\H�}�m�Wz%�CO��[	�@?S�"�w9m����GY���z0�,l��Oz^ZB@t�H�K&��y��d�\��W��7}����r��Q6R�*�Z_Wƙu=��\L�Y:Wӭە+����9D���j�,by��{�KM���]���h�)B��!Zvj�z���n$�C]�H��aFY����>K��&{]K���Le3�-dR$��,E^C�ՆcT>��X�ٱ�c�'4�+;ĺ��v�H C�I�H}v�j��u�&}��7қ�b����cϊ>N$T�	9]����\쵞��3'���4g����c��!�<���DcZ؝���@��*P���h���M͒��w>Y��Hch�/�Q>9? E* �pE<��A�ò`|�xTAr*�!y ?��1@I�2>W��c�v�|�a��ړW�R&�O��?��$U&��vR��R!��~f΁�ZδX,��d6j@�A,Z:��`��v&܍�A����a���sH^d6Z��-g*�'��7�䋲�[�qh�D����_d�(�h~�X�h9Y��NH�7���)�������mٵ� ��M!�Xd��NT$=#��0��vn��wfE�z�EvP5 �VMٙ�=�0�4oB��HJ aRg�K���{E���]7��Rǒ�k��&��,ROk�Q��j�g��`TfY�"��<�д�:�5A���\u�Qh�8��i�?�p�o�V��p�ǸZpJi
��c�؟�X_����,�\�o}��:\�S䈴,
 �]Al��I�P�my�Xf~�>�$A�"Т�#��Vǂ�w�P2�l�j��E8�@����1�����E��o��Ԥ�^E��:%~l�>d�]���ha�xЀ�~����pSݻ��sk�&Ӽ��sa�ilr����;]��ÌG5'��q��ٍ=m*�9�r���u~�����ѽ7����A�N�(�)6������˵�&_��ʵT2�5�>~��y�B����p�Gi/)�U�:���<�Щ%OJ�g���g��~�%_9�W��
E��~ !�=� �̾�~TJ]#��p�Ȫ�� bM�Q�B1�ϤV��m���z}�����(ęU��+��]>	�G���*IJ\�Fc�-�>�:T u����JFf�/��Z�7�D]�U�w�Њ���;���)�<��x�4Q���U��'�������'B���rV�j��m����X���eF�1�]���*%,���!mV���A·�_�a��	�)�!��I��j
��&Xр�e�Xw���9o�?B��s�X
��������=�G�E���l�_�h�3���뵝>W	�< �u�w"���B�A@o䠝!�K��}�Qoj:
��Qzpd��N͝�a�9�C��dƊ�M�ꢄ�ة#Ja�h*�Q��<o��ܴheJf�˧����%T�%M��1u}� ȪKf��=��8C	����T'�&V���e��io�:V}��l���l�Z'��ۮaek�Y?�S}?�R�D�0�9��d#��^�k�Z֟jv����e�e�ɣA�_�\U2i{K�c co���Rѥ���%��*�lY�����:Q�������C[շK���@�#g$��.����7�ȼ�Y,Շ����Z�$H�o�D��7�#��B��Ϟ>�ެ�r��ٿ��͹j��]w�����yB!cBy�'�X��PS0uN�ӊI�T�����؜߆���{�������LtS䐚��������`VL��@ ��E�1��@�0��~IR5�n�:�x��A�����M8(�� s@{A:,q��_��l�y퓟RM���M��>^"t�t2S �ۨ���>�����,bL����"�������ydݼϝ��nWh`���~�֙m�4�+1 �O�"��!�'PW������*�`�Iu|�4���qФ�5�z������h��qN;���af��J`�,��[AW��`�i�c�6�#�0Y'�I�0�)ӽ�W���x[6���J=̍�8�k�1�b�j�5^ǟ��%�P6~�^q
��ʊ��l	L�:���~�0��x?찇,n�yW�O���G�@�lYS�aJ���3D�����0���:�>x�̙Da�:��Δ�,����Fwл�B��5`ǠnHL{4�DJ͛�,!˺Gاp�mg��Ǟ�Ch	�S�/��Φd�֒�ë
/A��� ��x�`e��l������9�������A��%�Fkt+���P�v���f�9L,R�:�( ����B��F�%�2bL�8E���|!�:~���J[����G�'�Ƣ#ƕF��rk�F�
�j�q� ;2C>��$�C�9K���1�����V� t�I��4ii��� �C(J�҇,W&��҂�\3n�<����S���=�;-��?Zǝ2�P�?τ\:������y�d��2�H�MR��dY��_*��_��vfԒֻ��`�O��X=7����d���J��c"�tVD暟��Ԫ�L�����Mz�`񖪢E�QG�ٝ1�qi|uO�Z	����:�^D��Sq��}Vf����O{�s�vLq��q�f��R������M����C�O4(u�ێ����0����͹N��u�+��6!4��F�S>�u�����:�p��Q1{MA�j�@Si��c+Io�蕘D�������]���@���:3�\?�����5aھ=�?	 ly����lxn��˞�S�t���k-�)ir�Y�5@۪��&�R��ݯ�q�PV+~x{�܆�d���gCYnª�Τy3f|�D�Zy��b���z��_�����D�s�⭤�so��X5Q���O$����S� �^���ԀT�T�|���LJ�Ywg�j䮛3�F���U�-\�_]��ڵVa);>�����_��0�΁e���}�y��Ik�z��o�&p싎"����oF^�ia)����O�gz�Q ��>��&�ee&�k�n��H��H��[���]�K�zjr �"�3N�	tzd,���6�4X�9L)��|��3��tYu��V��?ɽ�-
�?_����wUq[k8�\H���	��qD��ǣ1{Q�V\~p7�r������I��C�U<�/!.�Ӳ]��tuW78��@�N�-^X6���P�� ��ҳ��t�<!�;g=�5k�?���� @��	�)w�OQ b7V�L\e�52j�,C����똍�������,�Z?$9�7fE��<�a���t_T�=�
5�VY�/�dOC���m�"<��E����+圍C��W�":{
y8�tRޗs!�eJ�x�BN�Cp���Ԡ����k�5�D����%�v�\Z2�l�} �^7���������as�/�W��,�5`8P�1Q~��6���̕(^���2�(��,\������Ai��ވ�
di I��U�p)=�S��ӆ���C�T/'~E�.��8���8� �T%�^e47��y��-���E�
P��¢�ʄ���)x���_@p�Nb����<q2w=��p��o�rlKSԖ�:ӝ4LʘcM���T��J������y���m�7f��m#��nkk	���y��dŐ?"n�#aQ,:5ź �b�Ҥ2���^���w���`��z`Ky����5�B���'�Y	7�,�uX(Ug������{ nRR@![Kכ���!y�ؘY��n�����L�L�"�~�V;��1M9�}b_��=>�<V�Oxn?CV�Ļ�pwD���n��P�گE��ȫZ�^.�{´�u��%�v�6]�t�і���Qc�b.��	΀	˃:�x��+,��Tj���I>������u �P����
.���Q~�ӆZЮ���:�V	Ɵ��e���H#O?����̗��Y�̩���ix�.t��93&Dw�v4^=��3s}�ѠO�`#3�I���������#��9�����}��et���5�~-�:��ܢ��|.��ja7�����	��k��S��Y��'��!Q	S8���sd�,��d��_���Y�SlX�uY��Y�#/j����mn�+<X[";7�D����V]����~܆�
��SS��D�r�r�D@�>,YD���^��os)�	�Ћ�]��ñP�A�؂;�N۪܉�./���]�|�'��x=�ƫ.����1��%���S��$�D�B�Q�a�erj]�p�t��#�4�0%�k\�.�`�|��ɒ�fxu�W��q:�5�.�b��������f>����	��F(��W��;8bwSB=�+*3����Bq��}dO�-y���xUy����M�`t�����������v�V��[/<���qp{6JR YO	�-?��ɳ"���SiJ�R'�O{��;tQ�PΥZO��`O;]�N��C�q�@��Z.W{l��#^��F>eE���,��R��W����3���x������y깸�y�m�� �b�D����W�D�,d�Q��DcY�Q���ī��Oh�x1�����nOE%�.�¡���l��А��{��_Ub����Q<}�@�р�/�^V�b� ����ؗ�^$�=����S�n���ENlp�>:EM�\��W�����p+н��[�ju2�FL?��~2���W�C5,bJד�`�L��J|lvΛ�Lo��y��K�wX������00�Ӑ$��8e���iC�v�����w"��D��R5�߲1 jr�����c^:��߮����'
O�s�\R�����	�M�����Ƌ�eʅ��]u�
�k�p>e�P���$�#Wr���T�<�Rz���[0�X�� ���[@�o� �K�)$c~�C������S����u�w�x�ߓ3^Ε"��w?_�p+S3i�x�P@�0rJ$��ª�)�>�Ҟ��y�������n/�̰�ٌ�]� 	�("L��H�|��|�f����V�JUc�t��jGizŢ�Nד�fq�����<:��׶q#[���Ͳd�u��뷥���ٯH�K� Y��2�pB�l�R�޳��iJ��ڹ��'DSK��[f�<�p�� 2�k���'+$#{�w�S�<�>�P�c h��*���;rKJ2�,6�k�Y`&Ys�bp9�&��؞a�@��i9T��_E��$N�G���`U�&xC��az��|M�>c`|il�9������|�� oL+0~�g�@��S��{�]#���X�˻��N�`�g$�]���zP��^֐u��M%N����w��m&�Ih��H��S!#�dVEY.m�`�ݬ�����y��QK��Ti����M��Y�(�̎��ܷ�����[{�8OG�P�߲�p�K��f���E��%���1u��,�Y�0ȗ�)��r�=3�,���<>䡀0U����x{��TV���R4*�D�L�a�]���k��iz�B���HoS���s*p.�Gn6���
�p)�K?5v6*z�~Z}��O�뇩���u=�ذ�mHZJf҉V���C�8N�BB+5�~��Y��6`)���}�[�F)�KY�ugm9C J9�Ѯ ��B����v��t^_=7�g�VG -6ݟM�]'���ک��c��gO	�),m!ɶ�H���Dޯ� ���ac3�#jHݳ���e�z
�!~`R:�Z�1&��u�i� ���DF(�D`fBΑR������W�"�H�`�H	<�(��V��|��«K{��<-�On�Ncv̲10�d�Z��C�B�])�sP�{�p(�c��ۈI��_s���o�9��z�:�����	�
��O�,�T*��s���8�<n�θ�@����K��Gό�vz�3!N(�Uo���-V�Y
��U�׏#z��Ĺ;�[�󰙠�LZ��p5��sV��_��}��L�2�)�b�.�1
����8�]�w���ݿt^��+�H޻�s6ipZG/3b�~�5m߽�o֣\'M~C/�2��+��8�Wf�hP,�	m/I���,;�n���SY�)�ki���>���~�Fjr�n�9�r�٢vnW��'݆�<�� y��jZ������%�	V#�����78�B�U5�_x��%dZp_`݆�~��1d5E���6�) ��MV���Ee�7�QhCgX��9��D��Zg�\�f�3���"GB��bD�����~����"��O��(��}'�����yF�W6��6�7��jk:���a6�q�+w��#=mV<s�w��k��#P�./~f�z�U�� ��{O�+W�
<����'�4Y�i\{���X���8�zh��WcP�4�ҬUb�	�%�W�k����<޾�e<�K�}��(�7]?�E���%�U���n?k�h�ɰ��֓�e'oGe�=:�NB��=P�ǐ���z��4��7��M�C%��$r*F�2��E[pR�0��z�#ǅm�P�+?�����]
��'�\~��7&�Y��f��[K1'����d���孉Έy+[��E	��v7�ɓ� ۸Tat���x:����$�z�+�/��D�����#�i���N8#��|P$K	=b�k�!�jǞUt.��[�&����4��Z��fr檳*��m1�M@�v!+dlmzWҏ���.aiC�$h(���4�ޙJ�T�X\0��)�C�\+�J/�W3F=�?��%h�|R���Z�T�!�!��*��=L�g�o]=�-[�7�ף��J\j��z��9�q�>��f:��
|�tVS	�h}Y?��A|[���9��W�+�w�N�!�`�JǍ�T�xu�s�쉆����T2J�����e��r���r�iu�	 ���û�JZ��-|�4�"���ȷě����(ٰ�g|����!� \A�{��S$g��-��ud��I�-TnT����)�?���Z�.a�-@P�"���*�^>����� �������.����oDd�/�WK��c�@�d���[������P좢13��aa�̬��j�rUK��i�����]�b}׉-\����+[�y�-qh��en�Z�D84����A���cjG�W�m��v䤲-��7�	����5��zVZ�~�!�jjy�a~�n[=T�u����-��E;���� �p���]�ɻ�)8F)�d��g�A��"�@���@2��-�"n�����ycE�j�Aɼ"��u6?�tέ&k�i�v(�u����]����^��ɏY�0�m0℈*ۦ�;r�L��`�*��?�C�ˤxf�a�� ��y2�e�T�f��-A�=��-�!λ��g�r���|�S�{#��A��N@ݜ^L�~\�d�9�������9kV����E�Bn���"B8���r}�#M�� Ϝ��m!;6�ބP&gj%���Z@^�"n|� '��s!�kv��-�|�pE���S�
��f�	����5=~N���1�4�ۯ���F�O��S�b̒3&#b��1�_[�O��޴��'dm��?�w#ی�Ȅ�I
��yF+�k�,��lP��:`�*Z%=+M]��R�Fz��4!�[����\�@���K){�\�ϋ1{8=)_cɓң�/pP0����e�W1��J�>"� �&� �?.~���lqW�(��@����	��}yz|���KX].F� eȰn�
�gY}Z�N���/�-�{�<([ �BX�mf9�����6�b�WSx=G�G��'������B�.PRI&��@^G�����}�z��^��~�Y\*|���x�A�3z��zXy�8%E;�� ��&�e�nTi�d!x����!�9Y�S���rn�>)ke���P\����7��mx3YHk׈�����E匇�@���̓�x)ۍ&������X��Evm�����O�����>��(�`ae�-B����A��U�G�sq����|�_�A�Q�{�P�=FÎ���n{ �ߍ����V�-��*�����Ц&�y��ѷ�Ѻ���[L7��D�N��Z"E�"���ǯ�##�-����sG�������Uw.Վ���:�	A�4f�[[�;���YE��C.G9��R���ܷ#�꒐Q(�o%V>u�^nѨ��͗}��ۆ�Ci�+��1�ʵj��HwBZ̅œ�#��Pu��\t������F����ʪ�Nם�_��01���!&i����4W�g�L,��R��pJ���>@��M���i�=~�c�=k������� �I	c�z(G�v/ˡʨ�'�/Lt� �.�P�J��vԗ�����g���cp�z�A+�G�`j�B^5�qJ�#��c>�g�d���8w���f������t��������O(�08�{:�^��23�:��w�J��C�Ǿ��-��ANeE����A��O;��T���I��>8*�%���/��Tw�}h�&��|	�c�e����|�6t��4F�R��s�lJP�Ã�7�X�Zv{<�����`��FN�wb(B��S��ľ�:���}u_Q{�8�{+!lvMu8�C� ǹ��=et��d�3�'�A3l���)��.LƉ)c�m ����Jh-- ��v`+Q��!"Jk�၂m�ݖ�?�Y
rj���)���6�Y�<$n����s����M('��˜Ў,z1wcg��X����7�tA���t�� 2�gtG5s
�z$ӂ\�-5C���א��?,9\�99��g5g�\F8�W��y�VP�-�;K��0��e�����w�;�p���5	P;��Pn*���w]-�CΖ�V�BW8~KJжN&�����c�X����pI�)|<����6m�������6�Uf��4� X�������n��x'WS����f�`$��C��yϸ�`�4�D�O/�?���E7�j�W�ֲ����&tRZIu������	�2�(/�{�K\��׾�D�����a@_Ӱq�r�/sqӽ^k�e�F9��g0t4��0����*u���`mγ���^KkQ&_�B�
a{���R̈́�%m`/4��F��F����$�+�h�~��Z�Sѷ���)5��^M�����ۣ��7i;�:�c��p�J5�NV���Y�P��X-j�CK���8}n~�$_nC,2����n6�9$tuj21�!��˚�A-�����)R��cÈ}.w6�@���pO�*-}�[���h-;w�_$�	��~��[P��o/XludOswx�l |�� l�����}�k�)��^qIǵ5.T�2�������V���뼕cy�,=#r��s���Dբ��!�����-���	���`>�vB8CQ����q� ڻ���P���;���`!�BP�+���M�h]���<"Y����NޥmyN��[��)[(�)�D[;:
U����(�T/�z*�����~����#al������\$3
� �QR���G.��>gk�N�b���u�h<��l� �?]�Ě�'�8�����yO�Z���ǵ}k[H��������!��gxȑ�"����5߃�6�;`��V4Ǥ$�%�6�S(~1���ӹ�G�oXN#g2�34Rܚ�S����=��i�kcLB��~F�/��T5��`I�����s��p�W�)�4"�P���c~Hn�F_�����ڗ�'��j�>WEJÀVF�U�V~2l[/�O���އ51@�;-=�N�N_S�r5�����Jt���&6��*I��Z&��|�����sAY���Y|.�q*�%Af���kt�ATz|�ԣc�a�j���欴��/㎭zj���
���S���g�����Z�����X)p;�� ��+>j�hk��-ф�n~%5�(� �/:з��^7�V�(h��O��0��|\4��\O��t#"]�VёrIf�8� \����)�~r���^�V��߬<b�;���S��c
>=�4(jT��n��W��!����H5!I���;��a�弊L,>�5*-���^�f��3��E��V�wn����48V���j\����{|{�O���h�g�e���b��|��e�U3�Z�BX�����1��6ܲ�hd{ M79~}2���yi1\9 �'�d0���#� �ɔIݍ-��aodȪ�Q�͏����U��Hx}�sF��W�4�jp��A���PhG��T��@�K��Q���t�h��h�+s�K��I�k
����ħ�?#�ssh��6-�h��'E:'��mԖ Փ��x�2���]��3s�j��R�]t�q��k��̓
]d~|O��DI�&�ϒ�a��%�@�;o��d���	��a��UW��}�%��o�j��`���W�+G8�"0c�/©8F1,��?o�����[���$V�F�0��*F��N6��ɋ� ��;�埳���@P�<X�a�v�N��y�\�|�d�}�N�ZCv�
��7�ѝ��^�����\��H�j��U���W�8vm�R��^�a}MV�8�� ��*�n��+(��PdA���=/&m�pZT�y��@���,?�&o~)~��$��^ �	݆\��6v2Y3[|��I��`�ڏA��7O�K��]q	�iM���44Y�&۴����z.˕λv��ŴKY* E���bHA)���:*Ŵ�q|35�sJP�#��_���Z�/�\�FK���kI�n&u=�v���;���R���5��-S8ߔ����4^:�I�����N�!��F��k��&7����ޟ�̩���Ml���+TB�ٷ�����
/xL����펾	��5郇s��<�Q m]��[]�c.gq�3�šQ��3o�M"ՕhE��\��<��=��(-{�ޓ�ը�J�q�2���˯�;�����F�\p��aBr1���'c7�W��p�u��W��	+L(��\�b �����q�>ǖj(N@�^�z� ����">2\�l&ϊ,�V����q+��!26Y���~/|�:�ӝ¸x'� �{��1��m����2��r"5!!�"x�ȯ��y�\z.nn�"+�r�����c)k)��d�o5� ����ti�N������}:tR�p�]=!�/ES:+��Q��g��i"m�Ei��z��ˬ�������7������	�,��rI?�*�iƝ��%����a���� ��)��1b�v�X�/0R�F�;����N�K�ucs�&�ʞ���,t-�Po�S*�T������>�h'�y>+��{'.^S�Qx��
Yo�y`�۾}�3T�2����cy��� /!�����a���.�	��Tj"�d'PӖ "P�=�����_ڋ����N;p�CD�
ixR)l&]���ˇ9�q�]������ԇ4���?�a�zr�fP�>p�ޓb� �4�+���d�`lB�ё�fRqT#Z.7���=j_��J�Z�wj��}r���{Ag���p�tB�m�H@��3$���f����;շv`��}�n ]yn-y1n!n�tT�{6�� ]���=>�m��&S��xG�2HK6���ފ�ړ�o�e���4����7ia�H����	ALg��RĞ?���trA(�TV�KE�a�D�T5Y�̨U�a(�L.�л�����}�,�SH^��M�dr�J���Q��>�o5���T���y}�l���*��ev: ��]I��4�X�I��hP���-�3����I� ��a~�9�MkH�.f8�$Hݐ稝��#T� ��ih��j����t{����_S���	 �\�BN,�B�褑���g&�w֨֩9����J�^�<���7d8<�^E}�bka��E���M	�G�^1.��a�Rz�oY�C#w��gG50��-������+pAg�l/�0g����]�W9�S��������.͔\ۢg� �d	�) ^i�A��[��|���m��V�7�Q�ڃ�1x^eJV�Q��η(G��y�ʋ0a%ؓޯ�&��*fŌL�$�}d����}�/h�+���a�����8 _����������$���N��r�~=��������)%��sr����.(S��z)��J�!Az,9��c�Hv�����@��N	^�#�����}�_����>��hxﴒ-�{F6����Ƴ�؎_�Y�fc&l�`�懅�q}T}
��?��s���;U�yJc��qC4���X6/\?�.0\B.��7���#Ja3��iĒ�V�W�PQEyč����?
�V@�Z�_Pl^��p~���*[���n����|�pݨt��4dd�~�eg��
�����m���́������U\Jb0V!"0�E�?x���ǟ�/�)�ưTh1K?������A['@�,~A�i�3����� ��}I�y���&R���4g��*��2gƐv��b@{͵T�`�XZ���QxI���?1��~��)s�_�:�lʣ�g�g�ջ\h��t���A�f	�̙�ބn�jB���֛[��:@�oR��hܞmGfʃ�]Hl�c�S	 ����+Z��[����*�gK�L�[6$���۫&_��=� �Ck��,�g��q��Z����/k���n�$x�,�ˎ�yd6FұmR��z���T��(2��v��'�h;�\xD���+�M�뭊��5r�s!n�e�^�A�_|ʄ�Xd �J,E����ߤuN� ^��(���=|M�\�.���8�IƇ~y���(a�� �4��Ps҄�����p^)�V��=����a(p���&��K}��j?�wg�{,|�0���.k���V����C�r�[��E/�m�X��׬r�l^U�΂�L����ޝ�q�}�#�����V>s�����L�:M�/�'`u�|��2�����`|�>�]B����_6>����hw�:������ƶ�:�Hl� ��� �����z��Opq��;I���zE�1��UA��G\�yT�^��ڏ	acZq���88��ea�;�ѽ�d�[�H~K]6�8Bu6�V�h�=Q�K���B��٘do�R�3]��A����^u�4��S�vݐ�.;�]j�"W����x��L�H��vPf��|�
<�{�WhSjf��i���5/qZ7��5�	hBbbE�˟d�z5�'�K�YZ�!uy��T,͌�KG��p2�]�]K2-�F߰�皽xq�{L��� �R�b�S���f�}�&�`��2=P�O�Q:�gι�w��?	����j��s
k�p5�!�^4h�I �]���|ND��'��$���5T���ϟ�b�u?�8�(�b��/F"#uѹ��_"��	�Z��)��TKJIF���~_}��N����'�t���1�L����>Z�������xӶl�%���aG{��!ξ;}�`�&߂�����ؖ@�sPr*`���u��M~��8�C��8�� )[WW�ˁ����*:�;D������X�z]Fƅ;��pA*�^/_�����#sC?Az�	��)�m%�h�SɵiI��$��H����៣��	�g4Y7��ç�P>2 �0���s��lsnb�������B�Es��𦧗G��U+����u5��B�2����b��Ժ%r�!�=�M�/\r�j�h����&"�$�zsx�L��F�ݖ�S�mpq�[^��}�s�I�Mo <H"��°a!_o�f��Ā��rI��D=������R��&7;88ӵ�p����ğ��<(V�Mt>oq����M6����s��#��N�a"k��h�������z���.���ݳ� u���-�'���-%�LV�q5� � 0�`:�=/��c�?�3<���ÎKY�L�������£�ɺk:�ut�sK����Uin��#��ay�z�����2P��O�M��ҧ��'��g�[U�;[~{��6✈�����^�����[�ۆ�F��#�d<-�݆(�>���z�L�h:]cc�U�W.�s ���	�(��jX(~O�������L�vq���S�]YkvM=
������5�'_�Y����$j(=͙�=�'�y@��G����E��Nm^�H�>�iwkNt6&�X֒1�<�VO9��N(A6J6I/����
L�ڕ�lʵb�@�����?B`�6�k1b❷�l��ۛDu|2� s_2�ː�ͮ�#|3��.��I���=���
	t����.a��v�(��J�4|���A��t������`WJ�?4*�Z�T�Fq5�"�(��k�X�S�a���?�<��L��J����I\�/�j��'���S�}3Yq03�'�b�6�$�ԧ��r�����1ѹ_Zz9
1�����b��Ԙ�����r��z"�&%?�7�Z���Rd��x�#��B� �L�S�@�����m~�ס��1H���|�]|����J�q�*
�b��y��ۋm�����^N�5eC�	W��^Za�T�<��A�a�K/����Ѻk֗w7��O��u!MjA0�K�����d�f�#�Q����;n��gF?�F)�B�9R��TJ����͕螢//�|�a`���"��ײj� ~T8��)�y��pl��QEu�Rf��v_7
�L$�=9�&��i�θ'z^2 ރ�]��s��A�;�e�)lC��qȇ�<�7��\�|ǟ��q�ܽ������ŜA�}���Y��L�𲎯�>7�zw��0Ҍ�����j����Γ���5�Zv�Q��~�HF	���{�jB��;Xx���{���$�!���@�T�|���_(/��?ci/��]eU�Y�ɮg�X�Y+NC =��\�l�՗�o&�q}���s�;+��?V+̛r�/EC�0Rw����o����@�K͌H�q�Z�����;C������j��\�5���h}���4��t���럧�]����9l�n5\�.����Z����y���C��O�D[��߻��hjXƅ���z<�	����zΉ�@���0�c8�5f0i88�,�o���mn����$	�|*�Q�R�)�0)�ѕyoF��q$���Ӷ;E(N` �����͞��2ȃ����r��pzVè�#EM�-��c=�(y�Z�N�;�xn�yS\iS����]�������w[W�F�^������H���4r�P�k�-�E����Nn�X���wb�H	���#�]�����!�P�..7x�6.F~sU��/�jM�-���,3�26�[���K��G���i?����k�	����x)G�3����e��l�S%���>Fi.u�O>\L�g�6�0��ȦY����NZ�����o�l�٬�϶wʹ���Mk��t��4\OWC�H�L{L�Q�w�e+��(���l�h_@��t����h�x>SQ�;��a;�^��q�pA\�Q�A�����rK�w����h`x�Φj�	x:�WEt�v`��r���$� �}�VP?���(�\���L��%e6kg�H�k9�I%D]*����@���HJ�cs� ��U�;62�����@���)��� \��nV�+�u��� ������Vv�������"q2Ķ5������.�m�ȭPxw�o	qX
 W)�	�hn	�}�O�4��8ˀB����ϲ��������7l�����;~�z{9L��WͿ�wȑ�\��G�[pU�I������Xqy�[�\,�|��5\ڲ �`��W��L4��e�����rғ|6�adO��l;���D��_�x�˝jW�wAX�N����?֝ӄr�\�"x5�F,�y��JC5����Y?��b���S\��A_Dg�4ʎ:���N]m e�ѰS*�u�i��U�rTR�u�/��Uxʤ	�r��G�[HLGh������x#a<�� ��-{	��m�$����+��2:":�N�L�r"��:ˁYʦ���Q��:�$��!%P���M��5`\�N�=o?��!�B�j���R��2]��[�C{����ZOKU����?��+�#קI����GQV�/_d�j�������B �Oz�dV���2�i<;�
<�(��t�gR:o���;�w�(���}p��(��f� �'/捂�acDGv�_�*�r*$I�����L���0�Ó�A�Z�����jmJq�%��ثZE�/o/gK��(�%�W�$��Ϣֲ���J��k��v�C�aT"
G1���=�ƅ�����Ԃ�;#���� m��%(r�� ]��9k2��:�y�H(t��H!;�e����R�_�gI�����X�쩤��1�]1�,C�sg�g1����J�ǕIH����S4�e�]����ZI��f��\�D�nxz��)�C/�g����^�6�͛15fJ��M}op�ZS�eB���:z&�M�M����R�D�9LG�4��C��?U:^t:*��`�۲j�go�K��+�k�Ѻ���d9Q��^���U[:c�����5��ݜU�Ā
�@��c�ڢ}i��/�F���R��,nA&��)�q)�@@�vaÜ	�JcA3������s�-khi�O?��ƪ��^�:����h٩�
 ����
�d���~���C��;�[!������>K,Q�]꾺K�g��o��'S�����5��W��*��O��=s�3��{�*|���	p4�\>0޷׎�`O�	�=v��`�0~�8~�����}���y�7A���� Jy�Kp ���V��>\�������q
�5l�5;��,�d6��,����*h���(�ʵt�] ],�&�%A���Bj�k��"���vmW��Ǻ(b����ԲR/��A����{���;?�Vئ�s�S	8쩂T2��'9�b���Sm�S�֢��G���9и�@��h*(�ک�l)/9�.h,R����ڱӱA���(����e*!�{�mQǶK���N�~�=�g�k����K�Ii`�߾p`�B�I�\�� ]�.f�>2�9��y�$  H�.}���_�$�����;�nq�#vc�!�݇Z�%�{D��� ��U�TT��΍.sT�63@���l�E���>��`��c����	����nڍN>[�� N0�²�"��M:���d!HsV�k���t�S{�D������-ح�q4v�	*# �wt����TznB�Gb���-�Q��?����Z�8���)�K�4P_��r��'u��`P����e�1� ;����;k}z��92�vl�HP(��\��g��.j ���F��\���i9z��5��	s-��tϮlV��X��k /��Ry�:E��C�ğ!��[9.F!�e������$�
8��o�5�R�_�泖=2_�*)V���j5w�FT��WcE����q�Z��`�W�T���J9����R]&]>����|n������/�A�I�K��&󎦣�4���q?����~b�꯻��0L�,K#��ٜ���K�����[��H&�0�Ӗ�b,��ا���5!��|������O�c9�x���L�����>�ھ��}����h���}�$*b	A���G{�6�FV{p��k	���,�����GP٠?A��'~�˯G��)/A���0�MWg�.e���A��G>E<ߐ���V\�C꒗�z���S"����&s����Z 
�����k��p��1ӌX~ͩ?Y��ސ�P��#�������L��1���\gE�n���c��/� ǉ�";
7�	b�vq�o2�c��rN�f`��Bψ������Iɍ�2.��l��0b^�G�36�?��r�R��f���i�H��2ڵȩa~�<��$� g�����H-3�.N��u>.GG|8<���ִ�J�%�ygj�O�ɲ��P�>=����*��TT�����S�?��G�uΒ�<W�,4��Ewm��  ��
j-�y�?4�I��
�G����B9�h�8fP�% �y�ڞ�'���Yޯx$Z�6o�|di�%_P#��L��_���ۻ�� ��	Dj�+t�������'��-���9�:A
��πett�w�h8jǌB�>`.U�an2ϓ����4=�BZ������Ü�����.���)k�sE��*(�%�PDz}�����N���"��FC.�_��0
�;쪫�������a�L2��馉3g���P��g�y<�w��6%�t�sQ�hÀ �[�;B��"?Xh�U��SJ�<m����q
CK;f������l>��MC�u��2�L�Gn�rR9�"2_��_sV$`a�����)�{�c��~��rd�I)^��u�6��d�ϑ (�߭��4�My��.v���R#sق����ZnURc��Oo4j}���κU $��=`d�_t�P�W۶e(g��l(��Qw�fwR"Jߏ��ő�:Н�	l��T�4��A������]&��?{�����8��(�7��H*���U.}�t���>���.��d��y&o�V�Lvi�Q�"N7�@�]����s�}oA2����� (���9K���8+����W�3KK�5���ٓ��_g�Ub0�+�b��$O��󃣊b�'����őN�+�xZ\�vi��L����&��L7�C1q��x�@9%<ҋq�*�K���Yߑ�P�"^�h����A�;��r�0i嘐����	�q!������(��­����Ğ=l��Dq�J˭yfm5�$�h���ʆ��S2����o����g�Qp�!I��Ym5�:� �ǍIz����q����:1�dѧ���K6&�.&��� �����X�,p��G�|�;�3�:BeZɼTCm�T�LO�����1����Sr;K���&�'�g�Ϛ����)q��o��� �<n��)5>K��%��2W MG�ʅ�t�����l�Tِ�aA��j.x�1���{�R��Q5�=�N�%�8Qy���9qF��n꼬aM0�1�0@���e-�
f(OK�U���Z��`�\�h���R�ه��x��#ӕ��έ]��cþsYp5S4Ŝ��-b��bϜ.��� Im�;I7a�&jibk��;���$��KAVg��O�)�>��@ak�u�i�?�U�8zYQW��{v��/��Q�*`.����Z��+r�ɣ+%�5b�L����1K��}�f���1�n=�����ȣx2K�H�/u�y��p�H��C{ U�Pu-ґ7MC�E2>�T�a<d/;�.x!p���+A�����$�84m-���d���(A~lk�7W�7������1�������wc
1CaE�g�ՠ�=)��۴{�ró���:ĵ6���mN������7 �u�f�n5�����-���a��>�#_���TB��6��6����ʥǿ	-�],~�qM���ZI�d�I��W�HLԑbd$�O�	�0>��:�^�i^RH&T0�{�޳�r��z��|���x�����:�o_�%V���C���XB�Mځ���_������Aܖ��jg�"7�Ŀ�Z�e�(_Ay)���U�^�s)�k���\��TDfȄ9H���#m�@فQ�)�<��$��EgN@��Z��灝T��4WP�j�o�ȝ�����9������b���N��'O�!���=��g��F.;����!��p�Mξ�=#wD��~nf���;c>ub�%���&y Ga�[rmUUR/9�=e���n4��Bw�%�m��m�^N�q�X�SWM#*�%���KLO��@��tA��#Y�^���j�������j7.���Z/'3�(�P��C�[�3i!j�hM�^j����,$�ڰ�����E4V�J����W*�9�&��V�ؽ�3�pQe����v�g5��0}���B����s�H?lP�9��q��Z*}7�}g��.�I>P&S���)	�A��� SݝS13�����&�ws�J���"W)����U<f�)Y�l�yA���,�A��-��;�M_�����lO����1#[�洄ש��.����ҽ1|�Qe设��y�>	tw��UM9���tH��F��%���އ�΍_؜mï���U�z�G�-�-޿��Yv��F?N;rC�$9C���`!��^O���/��EE�G X�Kg��p�ޕ�׊Bb�W��_�ÿ����Ul|`��L�>��f҆X}^��C��S�(J����ux1�T1�\��߶���h}��p����nje��j"�XE�3'��BZ����P�1Ƌ����&ps��py�.�
Ũ�Ӽ�k#H��OC6k�OQ���v˨PW����%ҭWf��܁~K�	ܤ��h�>�9z%J�h�#a��::���d	�M��3��{�o�s(|M��?�'󏬺���Ò`�+�h$��^��\�� `Gi1]tb|m�/�+ñ.~S�,���V��i@������0@�����:����.��k~�s����Ŀk�HLz٩�)�?��'_�{^�ӧ�X�?!�5�Q��)���\�MC�S���q��%J��ܿݗM�fN�ѰR����Wn y2æ�iS���vO���u� ���@	&'���T���sH���JO��k�����Ν�|�NU[[�Ƨ�s��'\D 1=�����C
�(�/j������ ٖ_x脳9�&�������~�ͦ��:�V)����X�]j�.�?0�'�Q,:�;��/SP�)��ƙ�CSH�A�I�Љ[�m~��:E3�JR�9V�p�������������PR�QO���[�s�O�u����?S9���v��1�M����s�+� �7P��' j�]T�W�u�ޢ`;�f��OIn��x.�±�D����s���O���an'^�06'2�v���CV�8���;�MEM��U
���������1��4�^[���*�$cg��8�����q���fh�wh�Y�n
�W�@Wg F���L]��F D�һ���STw�;��A��I�3���SxQ+D~z 
����g+�y��t�c|�٥�僪��~8��R�u��n�/�UJ3\^Uf�`�;G���\��.�zk�EGs_�_?g�x{��}�$��b�7����d/.?R�bD�I���s ���<>c
�\�$�< P
�Y�v K!�?��������r�.���56�('s����֯iC��0�=�
c��"�[�Z_w�0�x�)^��W����K?T���a��� ��n}`���/ax���bk��}���r�]e�����W�����7hd.#�쇈~�gR��\�˃LqB�e�h�D�Zޡ�<p
�M�y�'@a��8��
���۳���\F�&�R-vd:t�J:\��"A��p�X��R.��EА ��lb�I��
R���Z���N��
���rU���IA��">���(�Si䫗�l`�l�����_B�o��R��JA^��2C7�Y�Ov>�m�O�n��u��S�բ ���W:
�D7����g<Ks�F�R�7Y���t� rT���%36s�>��:�����P�C)�ˇ���=�nL�K��o�*�MĭL����EE�+�um[S��n��>�.��*3�������o�e}�s�ɓޝ_�4������r4of4�FQ� �R��F�.%�L.)�V��\�;��@d62�(���p��$���g!��4��o��Z����_`����(��8Uy6�j�P8��(�g�"�?g$��5��u�e�n��ώ4X���:Ȃ V��(v������o����F9(o���8ݿ:�z�jq�5ԲOG+��HJEC��ي����9�W���ֈ�u���<V1b+w��]��Iž'�r��S�8��[�����ޘZnt+�,��5�b���u�� ���ڌ3���ʔUU���l��f��BO� �%w�>(]�d�LT�Н��Y�@�c����E�	\n]ݕ�[�hF�6)�
�6j�K�KP�Rd]�6���Q��C�/3<=�]��<.DӼ�5�JW���Dn�=q�?q���,0���~�<�˄�G�#`~���� ��-��w��b �G�UVoB�?��)\P�s/�5�#?y��7�P�䱸PG
P,35����JO����6S��X���b�۝�t���T�Y��3帄}^��H�|�S:K	����_�#�x��?�z�F�c�-��u�݆�U�u�b�"�ǐܳ�7� Sr�oٯ����M�#��_A���ՇJ�+�z�O���(PW@F\0�\w3x��Qu�e�����?N������1O�֞���d�'�����"�JE	T ��+N�q�?{�^e�+8�������I����
ۆS>�=���P��\��Ҕ�f����70�C���K3|�?/�pq��N��OX�Ʊ��/�K㍦Lj�RL�]6,������x0Y�~�0siUL9L��$��h�g�N�K��7����9@��.�h'ϕ�~f�~oh��o�a:#���	H<��
��}<���Rw���n��	K]�v����K@U�!a�㳓~�vV�	�| /�á��!5���M�H/x�p��X��Y󂓌�L����W���B�l?J��/��N�����xO���Sy/��\<'��J�X�y���`�=7���Q�����~������C}g�]�ʯ��Q|6�X˰Ȉ	��1RsU9ڂQ�1Y�i�kr�:@��?�Vt���ϥ�/��b��:�lL}�����߼�%�A�����L��P��7�ct�=���NsX-7蕁�(ő1.q���oc�1�b�S����t?P�r�����,��O�~":^k����Ӌl�G2����g4��� r(x�=�1:zi{o�A�9;�B�f�:mV�X��{B,;t�Ќ�@ ]a&���|�:�1�n�!ɤ��NT�@�q\�@-=,J�L�@AC�h%�J=?iȡ�pW�0#_��52z��Q���h��C�6�$��v���R�r��Hc�g�����<�����M���P�oE�a�#���dA�><�/����)l	�׊�^�	S؋?��N!@K�I��l�8�PC�d��?D���$����.��eE^�lF&�Bjv�g�V�%)�J�:n1����Ԑ�Y���tjON�S�۱y����;(�c-�V��8��JGI�l��+�lL}�����u3�;H�>:B:���n$��F��skz�۔��6�T�?�&Z=V^lQ��ˣ�:Jo�`��!�	���)�]��Z�8UH�g܉�5J"�T�;;�F�ox�����gEYkE�Hv�b�V�>ϗ��Jo�?��b|$�/--�K^� �T��U٫��>E.U�4=��z�bF��'��P�]"�����ߧ�3)o�\���_M,�)�:O!Q 잼V[�����&�k�=��?��5���f�AN��tW�w%�$������EڥBץ`fv,��U�̌Y����^f����J��o�X�C���ۑ-k��6��*��r�,Z뀼Y�	�������
�t!��A/��2�JY��F��>m6�jς���r]"��P�NH���p>��]�pbb;�p��p���t���T�y�x�[�.s�2"��G�� �~8]7�^���b��~��%3����{�4eY[eTj��F\�{5�������ӆY���nO���O)]�6�k��O��q�r#�݅������ ����b5�L�;@P`����n������{-�����~�қ�1My���4��ؙ�h��ޗ\�?XI�h��b�OZt*%��0�۱+�t���	o
���/O� i-.R
0��#"�|n4��bڴy����r�V'=���=Oo��`a�@}�(�h܆v����FUY*���hQ"
��o���}4���)<��iݣڛ��>6:�F$,�
��&Ĉ�o$N���J������>[��M��u�/���U���W�����p��bC4@xuX,��Z��;��=@5�Z�����5��;t��s��9<+�A(�n�~׼�wW�ڛ����G�6�zqL��'VN�B#ca�q�N�.�,�'�K&��Nj��j�����\�E=Z��~�����J��fVO��T��Ȝ������*7T/��h @��؉�� �10�~�3�j�G���w��;y�Y��Z����6��g-'W׹� ��0���h�CNvz'7�͍ʈ���|��;��b.r���N'�$m4����u���Ͱt2ڋ�󺰥��#�>X��0k��C��3��)����������g�ҘQ�2G�"`LZ\���:pC2�iO��K!J�J�
 �E�64}@�do=Hk�BQ�O\c��N�ê��a���cX��2�� X�a� �$��v�a>��k���u���g��W�+x���
[HM���%�뙂�r��-��a1�m�X�~�ևp I��-��jn�)y�4��
\e�*�ۊ�4{����Xp�����~� I\�O*�:��/y�T�^�.�ms���^ҟ�1U4������ە�	�m��o׻Tbo���S�����!�w��c�P�\k=��x��y������dض��h��6 呼e�#_z��=\q;?/���(��i�+b���l�s��Z9".�̊����ժ��S�l#�Zѕ�i�w:��G��C���6����N�t`ܽ,B.Lǲ�7�U�� rH	�VP���Z��b�Ȥ�^��_���f�عZ�6��(�¹���v�#���k���\|�[�����E)#gd�g�Aq��Qq_�	S���x@���ʋ�l$� +�u�;O��o��J�m5���*<.$5�q~#����ژ�IP���C�j���i���ܹ��0��T��������-MBo��4F�%v���vQ^PY�Jt�vzf�)�np{�f�1ϭ����T`������O����BZ��^{�|�, Z-a�$z# ��I1���Ԇ�lL+p��J�������n#�.�Ů��>F�=�����(S9�pnh׸��GH�Y�-��^D�>R�ON]�</�hv6]��V�#0mµ�6!Y����˞�e6̫��%`�����P��g�zY���V�Q0��3mԖ���(��	~oF����Ss���[�n(�7=�S�M��r�C���0�.��kT�q�O��г�G���u���C���Wp���^��6�rj�c��-椞��T����}�a�L`tl��?�p�?�j5шPi�x�z��jk��@LGm���Tia��Y$�1��� Y�q���$�m�Tz�Cͱ�:N��B"<�-���m甝�h��Xh��uB��J8�yR�3��R��$�����m��7!u�(b,XCՁ	�͗��^��e3j�������-�0�����Ǟ�
��U�G�b��OKww"�l��@Йv���Hlv3U�c�=�~�RR^ʾ����ni#WX6��Wd1�T.k�]Î����c�����O?�B&��:�i[!�](g[��&�'��{�>짏 9?��o��m ���%oBk�BٕǴ"�(�s˟g�46"rp$c/���}	�:�xl���)��$>G�!���3�� /�Ⱥx�&� ����.��U�:z�ݷ�f.n�������~���c���D-�e-��n}��+��<`'j�.��H��B�/�ߨ�%�Ľު�W ���&��AP�	�랆��H�v7tL�Wr�2W�6Ș���D3.i������k\>*�2u�K~�L��=)����Y��sY�޿,�%��*����r���{i���l�"����ZQ���7���x)�����f'MS;i�܈C$h�|����S�� �P�^m���t��r���~����P$w��h�`�a��~�e�7��(���P8�c)�I���}�
�PB��o:2F���4��o��HX�$��v:�a�J�U�f�Rc��Ny+�_r�mY�}�����짠�H(,)�]لx��D�l����G����*���7��y-Y�O�*�
�TCE;&��˘k�/�E���{
��Y^�P�ʼ8�/5#��������[������q���Rl�֎<��/YC%��B�s<�J��pFɀ,Fs�FVa����?9^�5Q�.��qs���J[@| f%�B�!
,Ooa�C�s��YЃ	�7TqH�a��
E�;p�]jå�M�k��QE!�4>$D�9����������䓹Q_j�=�ik���"en����k_-u{&�ق7�k#�9|���΃�cDL<�U�)�N���T����=����x���֖G����ۼ��~��{ͮG���Y�"����p�`�><��H�>g�#_۵?���j�ڦh����,0C���H���6F��t������./n5�6r�d��ϛ/crk13�/h��*��F�k��l-�8�Ħ a����ǃ�?U�K�m0SE��fy&�_N�E��n$�coD5�w��c�(⿀�M��d��x�Ь�X(̩Z�jw�4Ni̢���ЗN͂�������\��\U9�qmf|��pN�ʢA���^��h��O-�jkg�q�Ook��{�p�,=3��#)�J1������&"ȿ1��q���(���_�!�)���^� ��3���q��+��%��l�HH�=���,9$ˮ*��Zߴ��Umc앾<_S�?.�o(���=��s����dQ�u��v��}7�-!��q�KԬ��nIO�F�W�`��"R5�%)����|M�]]�K�� ٨A��a��.��@�<R���q;I�/����"׬�|{��DT����h+\���R�L�H܀I�g�2A3��k��b�.�M�����;Ln��5&� �t�������'�^�Pv�	I��9�~���I:���
p#́�r�S4g3�Ҳf���G>������+7'V.W�=�u�sa�) ��}�y>ϪqY��Y� ��a~C���4�2TW�}��<?�"���Z��$��[ f/?4T��sy�[�d�R���H� /����^��]Yx`�F�iHa�/fo���ר9��������ұ�`}E���p��#1h*J�;b��6����(��5j�Ø5�lG�3;l�0XU��5�TpV�u���(s\��0�EA��g��c�]>�3���0���x?��_��d����r��3K�|}���M�u;��ǌ���y�8�*�)MA�I׫�C��Ec�0�H�3`�K��㏪����7�3`�Y�m!5)9�n$�y�|z�'�^��{L'm�~��[�: �)D�E������kD�lp�dc���E{$���榒 }@Zg��0%��xr��22������^�U�g/��=�A�N��ڿC<�E��T�!� >̈́�ݼ`�$�rZğ��,~'~jb��%�
Ů���Xƣ �o�X�s��A��C�@�������ϥ&����{h!!��ֱh'�;'9���نK}�v�࿤K��^���H"6��Tn#F��m�bm�M�����}�-.HK����W���ꄎ�`C�>�&�Rz�[��4�P�Ĉ�N	���|�j�m'^,.۴%\��+b'do��m-/Z���.۞����|�/x����nm�~�����T�]#|9���x�nd�UJ>E�	��"�N��h]��� yYx�?��n8�iq7K���ӽ�o��)��N����a��lj֓ ���Be��*���#�����=�N�[f��3���_�H��/΢������N�&��8�������<�����]:G/��j�t�H.�y��������V���IƲ��84a`߽�˙G\�>�������H4w���[l�;���W#�������(��-�<�8�ņ��Q����_�<B�_����بʵ}U,�7,A���-��b���'V��R���6&��\��&0�m�!ox��6;Ԕ� =1��6P�@!00���{�	ʞ`|Tl�8�m�����h_c�m� �b{Z��?����z��D�{��ۆ����%��v�Zō����(Ex~lv+��W���
�Z)uG�� ����Z72��F����0(ɦ�A�\y5���y���X4y�;���C����i�	�|����<g���Mr�p�ȶ���:���㊀�ˋ�燳d!�Ǖt�h� ����%��x
W�6e�1,=)���bӰ��B�5��xO
�vm��Lt���~՞�E��B_�#1�;h|��/�O�[�@�^�#�pR�)'���_�fBR����J1�*�~4hL�_{~�KH�R�ݏ%�;
�Ｈ%��3�7H�p{꜀�&{��հ}�x�-zB�r�9P�S.3�nO����Mڳ:�'�.��Ēm)�OS�@M�O���;u"m`w�nf��}%��]v�5^$bۍ�,;�a�y�SN	����� �8�_��׹�uR0�A��|	�CLD�R��.m̟)~=��
��|sU[����KP�	�P� Z�T��8�$�&.r-�Q��o��ˀ�4����3	�:�		5&hv�J�������%QDeC
�`�t�j]#.7Z�ի?�
q��)T�rX3:_��P����"�[�,�$-�؋�l�
�����/%?��Q�N�=S�g�����^h�X"��$)sՔ@H�����v�.1������#�t��cߟ^��.���ÑF��F�3f'�!WO�|/4Cޔ�vUOoBC�B+���*h���!�R�J�7DT�J? �P�z���#0ꫤ�:������?�Q ��|z��������I�ɖ�c�(�#��H�X]$W觿)^p_x\���Ku1Y�hLR�0�H�>Ȍ�_�9���������	Ee� ���%�@�,rE;�s$~�5����n!q�S����  F��aF���-P�5_���f ��7�v��%���7��+n/Z+.�
��3���H�>�̼�dk�M��)���r�Z�V�����@����t3��Q�9Z��-a`p�����wg�������ߣ�k�"�I��2�%m*��޷��Z�"�0�X�1�lS'r)ͯ����Y��9�FR|~
s1��+���.�G~��q��G�zp�xE6�~gf�!W|+�;�2֍m���}�Vqu3���Vjj��昖TM"|Y�eǕ�\-�b�%܎��?�[v�7��Z�`h���!=����tn�&�q���_*��C���+d��E��� D�;��5����d���$�~Ef�]�l��)R��!w��A�IØ޴�S�[38�r��#J$�J�pe��`��.6����M���A���kM�6��cZD�-J�}��ɒ+\ƕd����CY��x�� ��u^v�rQ��h�y�~a��y�}"R �O��Q�s��; [%�ʽ�E�>�S�/e_Z�0~��17���N�$4����-šch��N��=���p���[صc��,��=��`)�H���m�*IQ?飠:�y��;�sӜTɠ�.�k3 8;e�coO*�Ⱥ����Z��j����V`�k�� ����M
���t�-Kr1��`B�Җ�BBb ��GS�C�G7�`]Ee�r���쿖\83h�5�h^ݥ������b�"Q�>cʨ�?�E���sw](��ҋ}:ַ��Lb.|���)I!���(�_kk�I%��Qݬr��X.\�C�76�.�ż8�Cfri��ಃO�ձ������7���y �o}��SchR�:X�\Gn���RC�U��7�Cvf���P;���R?Fy��k�wر SӲ�ZҸ���Ѕ
�X򙆙ˊDQ���U�u)�q�*�W	��7�w:��c�N����RD  )lbu�D��>[����	-�c�4m�I��!I���G��3w� ���<`�}�x��&���G=Q�4��8��2�u<|��:A�it�����@Ո+6U�-b��rgin�8T*�@0���IB@�J'�f�l{�� �Ҫ��i�-��[dˣI8^�"�ٜ�6:�����G�oZ�۬���X�/{M��a6�&z��,��>��M�<u�U��{��9��GM�.��NVI*c���X�4��5��zrHm'6�m��ge��D�S�/'��;��cLs�p8U��4����.r�c�i9�P�Q;��N�Ih�=0b䂕՗6���O�(�s2��1ɡÀ���+���r�Z���9�Y ���2�Ҵ`߉�:�Z˔��-l���'�O��|.\�� �o�H(� QNR���Y�tfۜt��^4�\HO�<���u�^(�nx��\+Xp`����͊�F�l/Q|�����fX�w�R��()Ė���VȢY����.�� �'�R�:-'̕�kXa}�TK۠��T�W�u�����f_m��zR���'k�z�d}����T��?!�p��u�Y��5듋� {`���)���� .�rp�y�BQ�ޗ~�s������Z����5 �F@g�h �9#Q#񡽆ط�,��q��eXt��i�ܜ����-?ǋ��Z�Mn�����h���-c9X�~��Dy�H"1WL���\p���eR�g����:���%f"�;��߰lG(��zy��{f�tF
��M�XN��o:��N�ʗAܟ�oh}�F'[KT�~M�_���վ�0��23a���d�<=gN�֊�c��4=���P�n0�Jo��3�Ic1����s�7�
��x(�:����o�F��<�(%����o􂷤ƝB�s�B��N�v�k����������,�C�8g�l�W�˳�A� *�}D(��#a�l�A�l�PF��J�.V�y��>C:0�������ύ�פVj8��	�9���, a��a���7��U߄-�L�,������cZ-�F���<��G����z������ۙ����xn�8����6u�%޴�a��w���=�_a��?-;���8�߮4�)RM�%Ͼ1�W��ވxBt��^
Y���F���Q�����B���͔�X������+�=Vp��F���}>�&x�ÜpQ�Mg?/I:��v���ĭ[�V9��/�F�C���lcFrRO�nsX����}p�0m���<���1fuQ�^�:�|��0co�Sm�Fz�Xh�� ��!~k�Z���W�&�=��/��"������>o0�.�F��c��d��C�[D͗��e�0����g�LO�i�
g�̓��� .'��@L���;}�a�.�sI���T0�v�i@�@	����\�WX�T���okb���<�.\�߿o�����q#Hx�ϝ��F�zt7����O{�^��Wк�6w���G�r�ML�}��"����K��n|.23chޭmn�/D\����@�k��sA�^;���ٵ�"��e�oGT�%3Z�%mq�ֆ�C�y8b\!*GT3�c6rӌ?��J�B�\�	���ҵ��O����X��W?b�Q��[��ل4r�Ɖ���}�5!u+��K�Tq	'Ӡg T�dvgy�i."A3D��W̞�e�fUr�fyR�y4�Ł��k��V|×��׸�>�5���s��h6����%�{_t?(�|5C�*���}�@3�Xz�,=d߯������|.+�� �>������4�T�Ƀ��M�����l�0q|'1a;?WZ�by���w�	�^Fu��fMȜW�N8�[�l�?m}�Gn+u��nK����ȮM�"'�9��M��0e�6�Ulf��	�����*Ǘ�vIC�b��4�6ϓI�gd?���{�)�!�'?ۖ����D������(�g��A@��F ��LS��.�yo�u��o>��~�E�<N��S���F�;,8�%���w�z��������B\X��H��Je�|B�<�����)���r�g5�Y�Ak, �������Z��=5��(\����|x,���@��z��(Ճ�	^5�8��۹"��Awg�q���Y�=VGv�̠�/�!l�-c��B%������mW��p�cr.�ԋy�8�s��%=ޣ#T�e�8��*�l�:S��_;ݔ�L��2� ]"刔����QE�G��π�<�ؓ��7�:o���ؓ�88�q�=|���v� #�Dl�Ҷ�� ̠�wV �I�&�(�l;��!��!ά�NC�O�I�0��wJ���e��h�E�F����K i�H	�)�����!m�/&��98H���_p���~��exŨ x�}c��0	�Ч[��]�&HLr�tF �<����pa��4(?B�ʚ���2pk+f��Y��|��3���,�[2B��R����F�Q_J=Ŕk��(�%� �)�y6�6���ZS1��'1�$�u�%	�W�c�������)�%7B�gγ�*?����A���U�y��L�۸��-��V�9
����?Ҧ 8�-�u��ݴ�L�8���~����\�R�N>S��l�2\jߋ��ݯ �����&��陈���a9՝'W�����)���jh0Й$U�[���Π\��m5d!�N����gZ�*̕��G�FW�q�,eY��7c�FP�؇۰V~�����>o܏����Oe'�%���p�H��N���yd[�xyg���GM��7�aM#��z���X��F�l�V�[�Ӫ��ޚKO�We.}Ʃ}���A���?pM �����{�sx�+x����f�����ZŃ��;'��
��=%�'��[;�B�VqoCǲ���g�{S��,Pg�o���4�c?���G�&�q>�8��Oӝ�NG6��_Ihwh�~��vud(��2Ez���Bz!���������ZB�_6���u�VZ���q�����_��[ْ?�;T�W�N��
���#-��So���xC�5������&��]T1=s�D��`��-k���!b`�3�ѨpQIb%!n�]Z.�4O���_���+�J�¥��/�bۥ�M>{=j�a�V����n����8�o7��z^��A@��Cz����P�qW�{�:ESy	�������GU�3,�h%�k-J`X�K��Zz����-\��z�ڢsr���n�U4) ����2voIaժ�8�ְ��,�}�l"oR�tF��=��~}G��ң.�J0��2�d$ V4$��!t3�|�ɍ���ꩿ1��8��������e�h�;�sגH,��Ip�z���BN�W�|+����_�v)�65�h�	��l���`��(��-A����7Bes��G�>?m�vg�49�1�OSu�^�_���h�/��Q��
2$e��sNt��F�۷�;;�p@B����eC��SW��-�u�UzY�C�ڒt�� 5� �#?���LU�&(��bA��:�K�+I��M���j,g�G��z��/�u;xX&�����}�9��q�������4�Po�.��|�tu��X��D�7���2��N3mR�VH���j�Ĭ���NyT��Yp@�*��HF�>F.2����2�����ٲ��cs�	��.���9�t��sE1��)n{� ���I��ȱ�7���7��r�f]6���%�j�b��jP��:S��`�H�%��ӁyE	.��X��r��e�>[�T{�ܕE��@�gvy�#Z@B�h/��fjru���-}��#P��)c ��U���e�e}F˹PJa(�3���-���m^2�����e���B��	��_��m�5^�� �n�ӑ�f�@AF ��fA]@��������U���|�G��ݿ����u�F���D ��['n7"9�6Q����{�]�z��F�4�����=a��K2kb1H(;\�R�2ل`E"l�H�|k�O�~�n��P�.�����?�H�z�Xt9�`m�_&D���ӫ}ف� ��,���"����uy�Y(�+ٝ��7iC��^,�c�r��Q���o�T�|�H�۩w��ӍݓºL�mz(zf3�"�V����.><���j�I~'���%��[���o`w��4�z��B#�C�ODzd�-}
c�]�@΍%���� �ƶ\�$��+�9����|���u�~���C�l�&Q�� Y�,U���g�+z�bi��N8�� �����T���9A�m�,��%k�^G`2`*מ������7 ��	�Hg��[q��7 �K����s��k/q�e�Ǜh�~�1i��L��Cy�F�;1��=�6q2 �V�x�󸲔֛�=��ʳ�e���/�ϱ��x���Żuƭ�a��Q�<M�R��*������ĊK�j���̩S�;�2s�p7p��G T�h�4TR�k�< �s�\��`�����e{®\�,�����JJ#M4]���P�ǂ�Y����"B,c��إM��1�M��ʳ��P�w٧�K�x)q��}>��>�c�z�)J��;�fU/|��Ņ��X��C��@�+�g�ZBi���ϕP�uU����!���*��s3����9̻ߖ�8L�`��Js%�*�F��
ǫZ��v_jK�=���a��S`44'�@x�Ԕ�`��[v�^��(`i������B��I�E4M6�L�Z,p�fc�W�g����)��Ud�)�7��a�^$���t�Ey�@�(.���[&��u�l@���"xJ����\g![�&5��Ϊ���B�q��!��oֽ�b������PGJ���E���H�z�z�w�|Kl9IZ��v����w�gw>����:+�5��RC�T�2��8����6�R�ΤI�xX
S&��'X�H��I�C!IN��X�ne7L��K�]~����0�*8bE�&���gh4��U;#�#�8q����M��C �u���������[eog����6&��QjK�Rc�y�
.$�}���g#��gy?�(z�F�SD^�{�5�m���t��mu�/IM��х���������|h74�#;p^�>|@�/o��k� �P��\X�d��8I'�»�kc���c&�`�����,��U�9|��&��Iۍ�_S�&�����T�R���8���Ɨ�yj�\њ8�)����~�z8�Kh��z�`�A��
�߃����8��1��/1't"(d!ʰ,�_����7(jvmyl,M ŏ$Op,e�D�����MU�Z;�78�SF�2�$����y�qtɴ#�p��je�8�·`�������E5@o�7*��%)�%7C1�����#�Z�h�>�0j�i����!�rl)��纮't���')�c��j�!q�"b�'�����i���&|f��L袝���ϟ]��;B]s��R��x���g"o���2�\%E�|6
5"h$�����O�Pb'�O�T�4��T�����H L�I!��
{~t�f�8>�XZ���t����d�]�Ŷ4+F�Tr�=PL#�8o`��O�^�C� d�HO��s\:Dּ�,MԱ��������G����.�қ3G�:�(v�;L�Jl:�/�p�"��8.Z����UE	�z2�����i�T��	�N�E�(�X�!r&{\kBi��K�̥#V��SW�^��ې�+��]hB������'V�]ƺ0���6��D�g|��t؎/�Pڊo�=���vya�
�&"�=��w4dy%�|E�j�1G<\VzXEhs��'%��  (^��Y�P�`�{KR��>�6K�r5�����f�dc�5�Z�]�3�F~34<l�����Vԥ%�Y��q^���A�E���ӳ�N���C��ST�)��}
��=�ϟ%����Pf�e�G��,���$?�4����mQ<�/���@�6�oI �{��H��Z��3�o��c��:�<�`w&D�&�U��>�a�+��HSv]�Pl~n�<�B�����ܲ�]1(����#��c�]u@j�ԙD���1f�,E8�%&D���y��p���ǫ=9|U�D��U]����}�Q�h��]�~��� Ep|��iYZ�F����J��<�R�J�!zI?����rVT��ʪ��g��$oi����H�M�$^�4�d�����uƲ�sE}�O:L�ZC�Q�w U�`�5��?�f�Xq�����S��~�#� � Dn3nme��Ã�XB�^l优�.�d��G�����{{�V't�����4j�9��-���]��! ��(XZ�=����4۽0�p��J���3hj�a����l�_F�0P�6T�����NnHs���#�M��N�WЛ����@Q�m�ګ����X���x��xyF|�ϪWnu�hȯOAC����,��9 ����߃������8j�G���g�ߔ�c-j4z�ћ,EK���f;�Oo���&�F�Ԯ��4����� ���F��NPG( ������o��>�O��&`` ��~��;�M�5a3X�-��}.</��T_������9VX2���+�5D�*����+5�	�,�V��q��&���_9��<�O�W���߽x�.`�lX]��EyA{���17R*f���%�%%x�x��+ ������_=78z��2o�X�;���+`)��< ��̔��7�^,싶d��a1.�P��ē9{�2�̹@�Dg�]7K4���0����JS�J�[���t,(�2�=��̞�l��(��ݒ~�B�*����J�{tg�
p`���ONsrXBiK�r�݊�]�j_G�Jx�
q��n���T�G����^�8G�G�Ǭ��|i���`m�h@��d`c��n���8Pm�#��_س�v� ��7�槍뢶�s����(�~Rzp�A�@���X��Q,���P��*���j9����>���*c(���#��M�?i�O [��M�;����uSu~\ϼ�nk�F�+�`(G�H�k^����새�H�)���
f�^���A�����@_�������A�/������F��n�f`�b�:Q|����/ݷ�5���/�e�dP
�'O�ljI�v?�'jB�v/|��\{�E�/���&Zi�SN��*�T>�pք�V�������"�O:j�S�W�*���d���$���,ӴC��~
R��0��>�}��	���l[A�tx��0z�q����L���&ֱ���<l��Q�H:�9�$���u����p�
�P�z8�+�=�%<8z��FO2E �^������R�ccg!���/��!xpj��[+������$��W�m�B�C�z���b�UV�{��
��3�BQs�wƎ�o����jM�!�v��Av�L ."�A�w����G����N#�����ʐ �97�����NY�'dg7��	2��D�����'��<=8���%�����+�K/�a�zU,.X�C�X��*�n\o{G�Ѕ��cدC��/�+��IyΕ�>���u�C�d�V�O�����A��I[�޽8�W��R�^�xH�<�̀����0�^V�唃D�,dvB�E�*Ɏ`#E����vJ��q����/�ե�邐J �S�5^,2��V8�V�����i3s�i�?�a ���x�4E=ݖ5��&A�M���.���O��zbH)��D	s����/��MC}[����GE$�1)�u^aD\�#$3�X���D�Q�#�_q�;��D�!�N�����򤙼�*��̏�2:��?VK���j�o��&���+��@�XTR8�d=����}Ygײi(��̳�9��@�¸��|�G��Q4^�r�Lz5ycT��P �e�Y���;�O�	��1I�>ؾ�Nj��E�v_E���E Fٶ��F:�v�#;���rⷫ�P��Lv(`�C��z(Ӈ��ߡIpY����r��nÓtT����o(t��h��|��r{^0|�V�ꂦElE��fI&o�h��J\z�<��e��z` �|߶Y.��`]!�BCS�y�W47�)'�eѩ�O軇��:�z@XN��	˻�"���y]��Ρ�f��+�k+]�3�].
���Scr1*j�9����=�K��ͫ���yBMǣ�K���>���ϲD%���ڛ���L�ɰpG	P-�!��T^1խ(�_��q���!&��!joсt����=�1�h�g�oC�h~m���(H<+��Cn2��W5�A'Z9P��ׅ(<����}�=��d]���W��q�p�?�F�A�%��p2ԙ�����>ߺl���>�Ղ|k;}<������O���*��S�G�b<�uB5Eko*[��wU8-����M�PIu�B�~+�Z�܂�nм��J�'��� ���V\�#bh]�=���8.|s�c��{��I��95L���!;?���0R��<e!�fr�����3�'�ò��J^ޖX[O���2�~�U ��+[l�k�L���>ט�c9�-O��5���mbS�_%�I��z�����,e1;�ǩ]�
eb�����`�o�{5�\�����k�r"�"� �&6����9)�8Q��,�f�f���e�[5�yxe����,n\w�{�S����ʉ�ķ�PiA#E�(��s�׋Y�' ��
�E��
,�� �㦏EL:g�@��IgNQ���6�AF\��'􋄙��u��'�&�M���e�_���)8WѩRg��d�)I���U\��8���(�ʞ@�tx��{�T_�e�՗�A��ΥY�} ��?��cͰ��R#��9�� g�������0rx-E��ʈБ��wh^I�G�Fi/l�B�0<c����L:�Cb[�q+�b�><�,\�Ξ$�g�Ἒe�?\�Zׁ�ޝ�TF.����x�;�G���ܾoӤ�C^��u�.���ꂿ�iop������ ���us��Ε�'y����w0��O�{�$�y8
J��G�|��&�G�Eٻ�ď��)8�/�X���84gC���Wː~���.C�z!�)������X�?M���\���dr�TO�ؾ ��6ԕN�x������=�T��M�q�6������cu�l���1&���xy�(L����$����6�&��Cn��X�ο�e��� {x{��*׫�8)`.+V�lj����H��db"���晫�*�p�4����Si`^sȸ ��ب�����
û�ԭV8nX�m�"�{�I/��U:D����a�/)d�l� /^0g0W(yͱ�N`K�-,+j��+O��6#�ufl_k
XBu�܃���_���/-�R��:B��-��OXɻ�y�éݡ3�B���F����h���1���Z�LƑ�Ө��� 2�� 0�ogh��:�	�Rgfgyy#'@T��"�`9�z?�����@�`q���F���j��H����X�P�jGtW��h �^mhrt��=d�����On�N#�ѧQ��lI�wN&���LHxY��"yv��VW/���B������7���-7���l+n���g���r()S�#��S*� /AJT��x���"U��aY�I_�
K")���P#^����k��zx�mmPOM������mN(�����["�䀺��)T_J"�"w�)�YO��^r�{1����ݏ�]C�!X�.07L\͟}�N����PFA�3P,�A��24˺��J����[�u�!	༂j�&6�ϑ��w�=���h>��S�W�
��q��U8H�ɛ*��%-1>��5��"N)9�����[�x�/^� 4y�\��Y昋��k.\"�(VU�	 �=�@��R�!<={�v�&2���~*Vlak�m܉0k"�wB��������뜉��L��L��=T+ �by��.UPBUn�/k�۫�z�m���4:�朄H��;!go��2�Ą����M�w5H2�.�|Hi�$���Qz�Tn�{����^$%=D�6T��i�� ��c�O��$�X=�s�洰�FWD��k���v�^e�j�:��MDs�nr�7+]��Va���B�_ó�ogb֤$K��.<�������Ј 	\�3���5��XM��x�DF����}�<�FV�4.�P���'1�nX'�k���������Y�lI��t�L�0Eb���-=fy��Z_ׁS\�"�E��ʵ��|tm(�8�7 �|s���?�o��A}: 9 ��������[�(���9,NJ��NN&2?cpr��l(���#^֗�(V��z�c�a����/�Š�nUj@p�l]�i�h��IU���oXa k.�V,)��[����3�,c�:�>��A���O�`'�?��Ǌ�I�_<�?r�0�k͐S�J�ur�ΔR��9�bhw���vݯ ��Q�a��Nl�Q���4����ЀxuI�n��`STh���E�`�q�z��L��jq>oYem�%OF�gI��S?߁Ր��l�[�IT����۝�(H�=�D��k+N�I�飧��[�0.�:�Fg.��'&]�2�w�u߰ɡK��;���S-���P��A�v��k�5K9\��ě�M�%ֶ���vb�Z�W�t�m'�;��Y�?���W�-��ʓ!�SГ/=K`W�#+�Ll�T��r�U���+XG���#ѳګ
U���Sq���S�	�K��}q/�+��7OgH�-��{��D˷,�MoC$c`
0F�4�V��nY����jj0�E#��?�10�+�� m���S_�!��\P�����
��j>�'	5ZG'��>'���X41�c��*1H##��J��P�[̜���+���\��+�+��o�.H�[e��.�H?N�mj<������y�U�B��Vp��{\�z�63S�u����d���Y���q��H+�Eͦ9�MsLh,"����.�u�:��
ys�Z����ή��$�e(m~��a�}'�3q<m�ٟf�����������U��-3ɦ�$	{�(��9��&e�7����DO�̓^����ɞ���@9{��3[3k(�|X1ĵS�����*��z~��@��?�� ��e�@~��,1�4V������0:p�g4��Y�r}�����ts�j�~�"X��#��J�g��r�64]�_dy��ǚ��k��:����u?��l�0�������ӯ��S��>�^�q�=k�
�+��GZN�P��ͮ����%�HZZ�5P�~�����}hg;@^�&Lj���l�������-�^	���:Q�ݝ�8�w<��fß��.���}���x'Lf�tTЅx%�G���O27҈F�U��	[�n�\�kn��H9p�l�U�;�=�SjW�N��@���8�X�b�/��TӺN֗�u��`������(@C�մbDD|��n��_���&��=����juY���}W}A��U���<hp�׋�e����3����3S+�`S��j�Sp��A��YwB�X�u�D&Ɍ�+���&����|��ߛU�,�n2'xљ���H�t;����H��7��������ک<���
/��c܂���(����z���ƕ_��W����\�F3�1i��:�Q*7�&�3t�i�a��O�C�TzM|F�l�w�f�	�W߫֨��Oϣ��
d||�"U�����]kU(Q�O���u���J�*7�m���:}���Fn5�n�u*�"`�v:zk�!�����!<���<	�R[�L���6l���؁_���(�L��@{aɏ�v؅�Vd�?�\��IDGp�La��G���ma���ߒ 0G"MQ�E(��5$DU�h�4�{>$�78c� ��ln��d���mx!�uqc�>6�X�ߑk4�n�I�خ���dW�g��2���*`�Z��E���z>L��'b��q��$K2x�s'4iই�i3��LSW�^��/��}���������e��h��u	��I���F&���ڍ��A�0ש�Ӻ4�t�{��7�P�#�eӆ�z��y�&�
�&�C�^KGƊѿ��i������`^w�EY��L�Dg�!Ge��˓��������<�E�
�l�F@��r�GV(�˄%Q�Ku9h<�k�,���)�t^��u��\ϡG���z�E�3���Ѳ��s��0/�5\��`߄�W#��\��.I'�5�u~Y��v�T�2tO���lK{V������ '9�)j�e*7�VI���4���� �U�|o�:�z�d�����'�͞!B��/ ݧw�q�M�]���ʥS��o��:\6�V2A؅Iv<V�a��d�=����^��v������ʅ: �6Z�9�����	��3񊺇�G���2b:a{Ak�m!��.Ib�������Y���|��e�L��� /~��r���*t]gs7嶲f
?+dM҃ )f�y�?�Nq0A�b�'"�-Gg�62�rF�(�>���i\�������AdH�6���
.�O���Q!	;�����vƇ����`�:E���䝖e��s�!ߥ���y�=�qs�	0�X*�=�1�,�fC�����	+s�0�����ښ}|w��+����l�W�ot9�u��q���k��p��2�����)�X`B�Q8U����#��7����ǭ��!4�a>�����n�a�O�p�����ݵ;�&-�A�0�������V�TP��@�	IF�%7"=d�Й?T��$7�6u�eE�˭MZu�����xUܱ?�`�k��B��ɳ��ޠ˂��D����Ԉ� �{�V�*��-yhsĭ�nN�����*�+P�nӐ�I�K�<j�����Y�/��!7'B.X��:jzxk�r���Z�`=���p��r}<K�J0"�r�ԁdlA40���(J),r�zO�\~n�]�t��)���j>�L6�Df0
��ڙ-_[�0K^���s�T�-�ih0*��0���)��)Gw���u���w ]�Zj����!���v�-�c���f`L�n�����%�g�ri�"̕��m���e�J8kzU���J����J�1�����|pl�����5׻-�I����#�{'G�h�e�f�L�� ��#&.��/P���ι��G���J�d�i}_`�t,��TP�	�P���#D,1TB8AM��rU���� �K��b��U}��-�)D��+�j��>͉П��$<n��_AU�29틤B��q��u�4~�+c���ʸ���\]�������2��с/2'*��M�d�ڄ<�֠B�?,ON�����)_~���m���!�t���̓.�f��]���џ�`��G�Im���`�ŀ+��1�p*V�?��E�V�ڗ���mӋ�s4z��N��',T�"�'�y�b���o7��u��8S_��>���P#�롪J���Q��
�{�S�{V:��?Z衵|�@����0EkؗP�R�w��OxS�3�G�omr�?ڦ_{�r�'@��t������zb�d{@���'��,HKK3���s#_�c�#:�ǵ��*�#���(d0���S�C��Z� ���G�UyM����Y���7h����֒�T<�0]�(�2�"yͺ^�%�9_� �;af��-�P:ק��.�X�m��p��� ��ޕ�4�c:R�r1�6�`ǵ�BRniXo��� ���i���Co��'���/C�"IE�p���D���^]!�L;RO�ۍ\}���$�39��I3w��Δ��k�5PA0�zk�Y�3�ՑqLL�w`�Ԥ�"���;�aj/�T�|U%d�����ƾ��0
_7�pŽ1=��V�nq4ct��	��@Ù: �S�'���`����oj<15�rh�@����:�6�"�W�^��Fz��1	��=Jy��l발�C��<�������EiF���ϙ��2�T��w���Y6?Or!rc/n�i���!�C:�6��|�aH `+����y&��<n�[6�Ms��dl*�����|5�u���Ei��!��>���&Q ��}���\��Ł�3>�`O�Sq�n�e޵��I�˟G����'1@��T欑��S���ʗ*�ū	�Ba��O��x(������!��%r��A��g�Z懁(���满4Anܵ��8�G�m~�-�('�ɑwJ4�N�y��L��q��Ahl����[CZ%��]�e��?5���M���� �>%��(��X�#���Y���K�
2�+'���ݮ}���:�Ȅ����Mpm�g܈�G�
�G�}��d\V�/�K;*`qz�$1��?�c�������k��� z��
��&'G9<0�TO�E�.?=$� ��z)��S~�7�U�(�͖<"GJ�R�4#�^��Ԑ;�ڝ�l�o[�XqE߯=���0XT<��~��S�)�iP�d�����$��.sN0QyK0�-�#K ������+�hh��)_b�%k��o�0���R�A�=7�*0���L�K��'C2/���(�e,l3��jj���7�ݰT�fO���q�r��%)S�fs#�g�@�k��m]|�ȫUݠ��� �����Cp�(�`g?9���Am�	3�*�""����ug�)� ���ˍ�I�/�zf�u���Â���Ջ����:��6��35usp����{~��o�EW�+'�v����Y'ns�Sy܊��[\�8�}��<�Ĝi@h`�H���M�;�ё/O؇0��,!�!�˺�A�:T�v�bWp;?���`�;�se�8^Q�6֍�*��в�^rkwmN�M��o�ړX�b!��HFBb}	�}�]x��66'BvS,�I�yO��6*X�H˞�+�7�F]A.��Fi��`�������� �C�KĘ@��_hPI��&���`����|���C�l�2�¾���1�>�w~�J
`�C���@h�s�La���W޴S��d #%\�IJ�A��lلy��N�7DW�:�;ߙ�_����l��� �������׉%)��NI��YdY�."-Cr��\�ʱ�;�7��[�n��/���;��x��t�%6ʀ�S��џ�L������~��S�{��@'�֞�9�x�ʮ[�$��������������vt��'�pnQǗ'��8(��K����KU�w��ły	p09�m�8:Z�������@XjY���@!��>}�na _�pkvi����k�ӕ�n17D��m���-�敃by�mS�w-�8��QG�~�իΕ(E���������QЇ!+ڰ��v�H4�>���N���5j���?������	��mC�,�7�
�&,��q��������R1U��Ȳ:�/@�jߙ ��ߥ-�+�%�B�KT��t:�T0�L��	}��i��TS���G�sЅ�{������ZyS	���Q�I�1�_&K�8�~�����>)�Nmc�:�Y�CS9&��SlI�ܺb� ����s�&������z�������Ѩd9�W4�{�Dԥ�rENf�C�KH�x�G�pu����7M�<�0���X��(��BzGq~�yN���f�z�r�2%OD!�Ql�Q�]����a��.(�-�P�m��������z���O�?�!hZ����a���=�&�@�;�n�\�{�y\Fy*B#�s���]�":E�e���!��@�9���Ɏ؄.���hs�=&��3�$ÈOL�w�
ϟ�_4�_N�",�+Q� ]�������	�4�^��*LkrXa_9"F�w�ۃ0���X��z���f���yl�3�i<�Ǩ����{$3z�ԭ������d�^`݅��2�L���ϗ���[�|�]t��dh1��e���EWC�F�80э�CW4��b+��a;5�gΖ�z�9��=���p�q���}�/D)��M���0
Xv`�{m���9OI�d��z�|��JUuy�R|�y&���(���D͈����Vnl��~쮾7
G�93��q����fg(�(���z�>��	!m��5���&i30uΌΖJY�x�I}
���f�����AG�2CWj��˫Yg-31儛:Z3��3�����P��,E��l�ّJ(y �E>��R�͜raG(^5X�9K��c�]�{�����So�@�(b8��i��~�N�?���?�;T=Ā�U�e	\�[Pgl��3��f���e�Ge;:TƘCsWG�¦��K����& �H�^2N+ԏ���"�=��2��5K2.b�C�~T^n�����+.:����%e�e�@�
X���֫���U���W
�yK���~'?g�nB�C��ym�\qz�4R������3��ySb����Yy�`I1�"�����٥=��4R�q2�mR)�t_�!Ar�}G=S�ڥl�7(�=	R�y��̞
7�;��Q�䋻�GzR�8�!�}�3��Tޏ:���'�����v���b��&>"F5bQ�B������43g<h����轱�� �8+�<���o<������֔8��_��
�u�G�	�i��/���3��7
um�io(S�x���pV�²�s㿩i��|#�x��즁�j�{�2���]F���b�:��Yi �"�|Kh-�������NQ;�ϴ{��2�5~�0�c��\�^Oy�F|�03����~1f��G��'X��w�Zh¢�fW;�S���6������:c���㻶Ǹ�d�8�cO���.��I�m�:\�l�ݴ���<.�D~d�G�OI�����dS��S+t���u�2�� ���4�s�8�Y$P[N�8sL��2癃9����'t�M�H���~�|��L	�Z����S:Q���s��cC���`��������4z��L�QZ�uiNkJ�.��Ñ���C���l(�.������d�\��O�]���{�����楲%_�!:�z$���`Z�h�:wf�Z}���.�?�/��u����Wᅅ!%ʺ�,�}Y7"o���}QЃ��/L�x���?Y�{�&�J�d�{S����Y���b�	c�2��r� z�f�򈒁���rӔb��r�2�u��H����g����k�Z���	���m �*UX�u럁�ɑ�����+4��0xg9�����C��M���;D���:%1�:�`�;�s#f"��@�K~�_���f6]�+��Ѷ�=2����vC���q�mG�2Dť4|�!���I6�?�v�6�]HC~تq��;_����D>8yk�ױ墫OB|���bd�8�Ӳ�F�Ù(��*��M��p��\���A@�,�Hl�>dX��7s�!���|P3�	n��C�xn������a�룇2��b�v�}�$Iʰ\J��oZ*O&; ����*pR��G	`"��6�_M����}<s�my�J[6p]�e裼Cz�"�CwP�ٓMFɷ!�.�PJ�uHzT)��V���-uA��q��X�5�[M��� �U�5�6�V1;��v�&����MXs��× ��~�{i[V�h�2,K��3�t��51��=u��>�L��e�S�8f�"�5����n����,@}g�\����s��������{o���o킙�6wh���(�WO(E�H�������Qhy�C���5�k$�f����p�i�/^L�EGi��\�\k��f=	��}�4�3�ج��UO|`��x��B��)�X�}8���ejC@�a���A�t�
���c}�O�.�� 5�9`R�n��������)�p �Ғ�8�P�����rGA{�s����GlYǵ��\|�#���C9�&��������|S�#v�4?��UK����z��;��)��0��Q����
9`�]�#()L��'�;�b����cä�)ʥS0B�˸�\`�&��F�J��{��N��x�ϊ�{~n� %�Tm�܍�W�i�2/����p�3�5�����~(��	�y��k�9"��S�N���U/��C��Bݸ�6o_��R��k��y�8���f\�/�$�՝�y�K
�����8	�	L��1HA�#������N�,5g�����R��������5�H��P.C��;E)Lh E�(�jؐ=|��������d���{�,&��Q=��G���j}2�7��T�"JO�t��\���|���y�2�-�z���탎��@��g�3��������&�(����� �Whk��/-�L��Ha��u�)�e�ʚ�N�$��A�!N@��p0�A�&�=���4��1M/���,�>G���aQ'����a��)�dz��&	���D�5R�����(�9߇꘶��Ng���,�h]���q�m:�0���7sD4���]��l��G��j�#�m�E|h*u�6n�Q����wq4x�&M�I�%I���&[@_����U�o���w��"$�*�n
���0<wlJ�éT#^Cp>��p3bL&�joN|�����)W���]j����L^ꪙ6m9��BY��f���2�0ڇc���y0�uZO��9�<�;��y1��Q��D�@�����<�J͛���GfJ����T� +9�JB&5/I��o-�J��&kL�Z���!���?6��Ѣ���<q8ʮ���4|��_�Fz�;+;I��3�.Z��K�t�5�-��_����M��$ρ�Q�qJ��@��b���>�����\�D�v�����Ԉ��ρVE�k���n�ƺ�����-y4�Aeé�
�\�kZl�,C�^O�	mDK�K�B�<�-C`ȝR���9������Zӄ���'D�!I�0ѽ���?Z։�PM�q�[M"׬-�X���~� ��x}��>'X�H��ڬ%��6d�"-oh���}�v�\=w�_%�
��<�Ý!M~S���#�:qa�>Ұ&�m�ZZD�a^�]Wg1�.9X�y��S�.a��c�}`Ί�7a#/%���ls�kA�`�`��Zlܑ�̀Z��*�-�)pQꂔ������7��,W���h�׮x��:g�V8
���ۅ�nY\���{3GG�9�*�Ռ1��O�����.3P�#�y3�_-��e�[��;%0R45�N��>�ϰ~���[>���
��t���F���Ww&�d���u�D5��<i]_z֧�KrI��O����W*\���F������kx���%���o�`�_H�Ϝ���;�:���!L�B��)z�0r�Y1�Q����W>�)�W�
�d݉عF��j���T���&��Y�U�d	ʠ0�<[�''�obU�dBC>�և�`�ڈc'���]0
�2`���;nu�o�Z�$������ɐX��"v�``���_�mr�e�}�q�9V-�GZ^�^�|��lO*96�)�E�k��,K�c�).�&ur#|�Ѫ�eҴs���$M\�ܔ���{br�IB��t��d���`/��Ur&`��� =�b�[H��2��e�U�`�<�wA��f-�=p�MBқh���7�3�xt����J�o6R��#�t������rzkc���8��?8���|tPӁ0]��M|B ޲�J3�썸���`����>^ݜ���g�_L��fv����B���0���n�xu?�w�Y�E ê1�d�<�}��@�h�oY��M,�d��w(m��|��3������˼�|�>�].b�TI�+�H��5e�<���,�΁{վg�Xv���I[ �u�P�������Q惁�zR_�
�T���$�%�ὗXj"�fm�Kh�/���x��T��$�T'GZ��xK�%{�u� ��U��K7gGt��G����N]�FK��4�5�f�8
�$���3��t�	M��[%���B�5���V�x��~Y.��.r �]��i���05����
ewB�_]��Q���:J���9.
��{��_�ܙ^��"�Jh�>���צ�Pq9�q���Y���0LK0�ˮ �'§��?,����ީ�Ċ2S�%�/�wU� a��� 2��1-aƒ�&�g��r.<�"��HH�U�kI���s�R����@W�H H!��GyX���%t�����
�(ؕn���(m���3�9%�P�լ�6�B����p�V�Y�rR<-��5Ccq����B��nt���tM�P3��o(a� >%�d~s��8a�+ز�h�β���}�9|f��eM�&C�+�Qס��a�*��yG������[�ZK���\���Yʺj+!Un����lI�j�y���K����㮞Sp��(I��79��Z����B�J��������z�Bk6����h1�2=:X􁠘���Q�R}���p-����uC-�w�4��H�f�������~e0❢	�����3�C��xdl���ʔ�kyH,��q*(�ہ�'�f9kY9�
�v���|՗H�JSܯi�Q1�-�x~�bu$���� ��H
zjM����b��n�����%/dc��iN�#���<��]�*�m)8!�}V�e�@�oE�[�����z�,�c\&��߲#����[
S�Ƽ'(�xG=���q��G�*���I���4Xv�R��n�I����Ɩ5�HQW��<��`._O��ީtu��'Ɵ�ݧ�"�2Pi"�-iE�����VX��v[�0�WD��o�ίP���e��6��֖��ߎ���nR`��I������ybTK�x�6�ӷC��"ė�@�7��>���J�R+?D��6�v�N"��u��� ��:� '=�\�+�e/8�!���-�lcx�r��A�q�pںT��Ǝ�MǏ�Ә�K
�����i�e;���.o�����NGA�",�rk0_:,6���k�V����߼Gӯi^D/i�r�b�Svr�����k�C��$���]F��;)D1�>���S֕�T��kMJ�����Gs���Ӱ^iՄ\sW:h1���;Qw1��Q�RŤ��Ʋ"'��0���ޒc��aʣ"��h��Vb��S�7`Y�@�T�;.��ϒL��1Ϥʕ扙S�x&I�E��)-�q�gw�Ƕ94o�SS�n�[�޶��i�`u5�=��d�LH�\��D���I�~�}����]��[@���;�>ؾ	�Ix�JMJ{άQ�v�n�'j����o�_8��Z)?d���C����" ���gN|"C��B�?��"�p����bl´��(�$�ٌ񤜰��TB�F����L����󄨘à~����L+7�8���CM+�/!�s��tV"jq�R�1+cX���VdsLAv�%޶�\��z<���~l@����n��>��=�E��M
h�1��1��{@����U�M�Ok��]T�},T��f%G�7lo/p���~���Vm��I���3hr�amI��u��7:_G�Y�l>>���b�Y��"��n����:}��
�et&�y��L�Iҧ^����6yqKl���H�m�;Ԍ�)�y���TSk�2��U1V5-�Q�;uu{W�ǩ�^���������4YRA��kxN�~��X�pۤ���:�˫e�m���g��XlgU��7z�J��������S.t�P����y%������o��|U<L��WW��|�z-_���,y�`-���M�����Q�R��<��]�n���b0��.�8�5 �Yu[>_yTix���E��{˘�.����8��+&iZ{uOo϶ڵ�����:4�6��؆��>�� MaA&y�ͺ���&
����f�ݴ$���1U�ر�žѡ��a�:�<Y"at�033M�9˺8��zS�٬쌕i��������>]��z'ax�&��5�_87�n���r��_��)3v}���3]u��5��������r6�*7<%��ۙ�����u	]wd4�A���k>�W���t�,���V��x^���g0=����m]��^��d_�!�GN!�����&K~��%T/��U)3t�IQ�I[��>PX�����0�����R^L_�� �YB@\�\�p\�i�"?�Jzzq2��~3W��&?L*1��7�1��)ow�S� ��-��TQ�`�u�4[1-��{0E�f�W�\������^�+��4Hf	�ޯ�;3�},����S�y���9��	�.�֡��է�M���\�C�@��b����9=u���ưZ$䯝R��.7a���wo���n��v�4|�y^;Z��o%5�[� 2�#���� f:��Y�A?�����}�������d |�շ�aWD��ZV�On�lx�1���/N�r[�"Aђ7+a�s�G��W�.�W Q%� �W�8��7�|�U�$z��.r�Bq����P���˻���F[2(zڶ�Ж��9?��;~�^M�Pb�g��y�ڽ�v<�1����w�Ə��ԑ�a�=فNC��1�ǁ���e��=�戧��F1���DU�q�a��Xa��`�;fD{@rљ��}�ه��g�CV.����(Bx��c���{P5-?�� έa�_8n�۽y\�yY���N���t�3�"Z���9NHCzƛ�k��IQyg���2E��R���j=]�_0���ݾsk��&����)���$^(��C�zZ��nX��ɭR`��$H�U��H�y�� -$�XHޞÃ!zf�D�8��}-q��Y�ͻ�mL��2A��rek�+��ߪ���*����x+�2�ʅ>�F`�9O�<]�i�KH�J����U�(��=%A��#4�y�h)�;��^��ϟ���Z��|��>����j�7�O5���r���;J�6!��K21b���H@�����
�BXQ�s��\�"�p����RRn��Wt�h�I���WI�y���;�p�cѸ,�V"�Ā���	�8�x#Zs7�D���>���� /��s�.Nk#d&}L�.��޹���u��1�C�N�3�M᳿n�;�d~+��͠�B1�!�����T���I4"ĝA�\x/VÌ��"n�l��=�͜~J9A���~[��@��*��wNA�Y��gs*��ق��L���B�"eg:����3U�G$�6��^�����;���ѱ޸jG���(б��&�6��-��	$x��З>�Z�J���s�&�}�g�6%4�n[����Z �!mI@>Vg)Sd>�WJ�l�Bz_'A��s�!���i�E��ߗ)��[�M/-�0�T�V ZV�r�v�����tQ����F�W��,*��j( 4+�(��͓�ϼ��|� O�x⎜�؂��ۨ'�?�^ԥvU�����(H�<{\�0�zw��vw�VӐ��0�>�/��Oj�g1�����z�!K���XѶb�"6=�����~
��g��8�B����Z������tb�Yr�#�l�ly��EIb$�-����L��ax��b/m�2]q���g@���o�<L�]�\�ʺ^�:��y��#�+l�"^y�@�����xL�b�;��~�8��=�����5��0������hU�_&��>��@�FPXB�����߮�0�x�� ���ƛ:5t�Sʼy��
��A5�4Bs�k�_y�$�d�˗�ѴW��'H����D"��s��+[a�8����8��\p{�F���Rn�CtZ1jo\Y�Z{�tbA|i�Z9�}�~�o��p��jy�@���=J�q�0�l�J;��: h`&�J6�F&���P���[Rg���-Day���,�k�B�){.��k��ދ+&���aۘ+�����#M�W�%[Ƿ�y�*�c:U�ඥZ��Ig!|@~�K�ps���Kh�y!Ҁ��;�^k(�
gwz*���)��j�;5��ϚQ��w��Ke�!�Dg!�	��ECͼ/�`,�Z�KzK8 ���p��ȇڷ7P8�(�Კ�mB-�X��C^+{�V���n��_�4>��M5#@\���Z�A�$S��'����@̱R��O�FK/ȳ�����w�R����l�6��}j����"���(V��%���O&��{��C��<Ƶ�hDto>�^I9'�U��sDUc3�2��$�L��������*;XI�!���碴,p�iŨ����1�l�\,%��]q�z�ĉ����a��u_Zֹ�o|&H���kSX/ �{^��V3�������e�T�Y����_�"S��=�{8+y�.�!��#�/�5���'��$d\Ƿ؏bԆo#�,���\�E7w�&ΓbQ�������
�����/���"�^%<��G0�<O�t�������ܖb�ɜxI�K�oV�͝����pٙК���l�u��찆e/����w��K��?���l�R$2��Ѽ�+���Q��lF��`x~ �1�V� �]�6�È�6*/2i��PZ�:��F��h���?��U�md**��Erqk.���D/���<xt'�ͪ��ň��9�q<��0�Ձ�����SZ%��4,�, �"���{�<�ǒ���E�i�n�ҧ��Az,i�O,��$+E�#�O�[g�%������y�NS �
��g��Ğ���.<�\�M��t�r��5(�E�8������9�5�t���#���"�h�ZY��o)�p�m�}ק�Xe;�zBt����ZmK�Zmg�Q1�_�I6_�.��X�+��N�gjg�Ы�H�W�m%	��NoV�4f�H�?�^���%�IOw����AU�T�M$$����O��Jpى���9e�{v�{O��DՁ��_�a���	�ޗ<3.��F��c���^��8=�8e!�������;S���eY�Qhw-�aY��d�(�w��2�%�6�WX~?�`_�������Mp3��><�8�Oί2��8)�D�U���?=���D�x���"�#��i$�Ļ�r�YFˑ��(�B�N��`k�)�n�����MU:δ�`"$h;���v
޽�7��'� v8�ws��g&9m@9 �&�7aygb����l���N7C���C��E�Q�-����x�#V	b����r5�L���e�&�6�H3�9��R�W�Z;���rO.4���c�}����]�3;!�����h���|�<�Ͽ�R�9����0�5o���>!Լ�KC�'�HE�}�N]5V/�����T7��҇_�{��hu�&���8z�xf���0_a�k�zK�^ m�R`��4��������x���1�v~�È��a�o��=��[�;H-�RHt���S�p���*�����w�b��0����v�ʉ	��}�����b5q�Z]�곷vJ��$������v�2�������e�q��H�h�_��,gr1��J6ۇ�ԅ���5݌S���g��g3��Ϸr"g��%eKZ�c��}�	���X�ˆ���ޠ)sn�	����B|���X����#����	�*�=^z���Q@f�fQA0�n����K�O����z��&2M�T�Z�u|�:]�JAM+3����O��CD�\mP"�Z�	�Q������R�"
�,O��-�R;ۑ2�^͗,�+�aUҀ4�St'U�,Z���W���� ��|�#y7Xph��U�&M���+7
U�C�SBX�f:Qib�_rN�H�p�
��+��m��1�0���JL��͕��X�9o��;>V+'�G�Po�
S��>�����z4�H�"fzGTjT���/?�Ҫ�{j�뽆�j-��gԻ?Y��c3�5Pz�6�$�{����(��{z�E����c7Z_G�!eXo?\����g&c/KK�e� ����l����0\ǘIGui���M"��y$���W�A/f|�uu��.}�J�f��U*�KG��ֲ�>,<�B1�Q �hc���+�S�b4<h�W�8n��t�|G{V{��xX<����밳Ks#,4L4����X�Q����}K˂J�^/�����wR����y� ��W� �}q�����g$إ���;�AɄ῭��b�Ys�#���N�3g�WDd��Sv��T^�T�m�Вa�]��9𱦠z��sm�X�1v�s��G�����d�r\x8���"�۠E��B�C�p4�19�1N�>Hͪ.Zf0�c�G�"�Dؙ4�^�oB�ӲL?�j�� J��ݒWI�H`�p����6�I�c������g�k�ĞG��Q�
ˈd�F�oB��"ֺ��V�����8B8��Ƹ�	1���s��Ol��t�܋����ΠMc<uc1��.���-�^b�&���>E��ݸ�H��"y�c
yIo��g��Zʻa�b�i]�nv�C=��ʀ3�* �$"����K���	8���W�ḷ��5���i,�=#j�
�{+ea��QM
F��5�����u�5�<8su�bR�}��K�_�z��#�  ����a�=�m:��sj��etIݗ0q�ꂈ�|���̪BD��`���Ü�p$�x�]��U�*y2lþU��}�3�1{U�����S<�:�7.�r�qhuP?�W�f^��V�~<z	H�ߓ���,M�㬧B�� �h�y���B����Z��-��n"+I"�r�<��� �۹D �b��BGq�~$UFκZ��w�&ϕJ�G��8Wg�<�#?m: �U ��v�A+D��ƝI�eWJS9u�9/��'V�
Z(T?�o�,T��U���U��BZ�m��{�M)�$*7:�5�#�u��J/�FAm�h�n�c[�b(rt$��t�M.�#����#]����h���o8��e|��x�A#�o�Y����x��B��5.wM�B��Y��������Hƾ+�
��聇�̶li $�j�+���H�#CheMv]�"�\wߤ�I(��x�.��74kNrS�R��o�߹�2�əi6\ >q]f�����(��m�bN�܏����B���w]����[9�}P(���ͯ����"��JV�B�X�Y�����5���,�$��e�{�vh�!�Rzk�z\()�,�w>ϪZ�$#Ů��T����_�F��s#��(�]~
H/��@>&!�k���.;s�ڷg����d��8��ک-4Q�\y�{�5�x��a���"6�k�+h<��z��QЀV���L6������S�����V6�`���C�`�0�4qHB^��@�Ķ' �����H�!M�Z�qXʄeO�X���0p����_�мVN�L���4\��Io�C�02|��G�Ͽ���G]�q�Rҳ����CM��gӻ�i�)��7����g�&R��<7�a�]ǻ"��8id;u۹3,6����C;{y��1�[h��Q ��(�@Q�	U����^����T��MPf.r<��7/Y��*	3�ׇ�%ee��W�(h7 O�k{jJ�j s����ot6UrOc�T�pĈ��Y�k�H�� AĠ4�_ZFn3tb�Ss8E��0U#�1���g}=��ƹՄ%��|�,9?��z�d�4G�/�GJ�%W�k���姈����s�w�iJ,�'k�dt������_�;�/M��k��Xx�����7+��Sؒ�jxlR�g��ӈ�1�Z�F�~G�兏�K������_�р��w��',�B���#�>�}
E�,d�L�
��S/D��/f.���t+R�*�S�<������|Y/��k�'��,��i�%�-g?�XR���G˗4�r˒@2b*O�QJ�1g����Y0�]g��piq�^�I#&	�
�F��O�F�@3r��4H�(�Z'�LCr��G��$3mo������K�7�_5ks!ZĴa�~�>��hCyrD��!d�i)��J6�b��k�������k�~�MYnꂪ�Bq{ ����t�^�6'� �wja��b��Bp��vD��@�) ��g4����R�pz
�!��0#��8��	O�Xa�"��#�\Б0�y+ �p��<�h���K�CK����"T�R���<ߗ>�q���[�P,�o%�՞,!yF~	�d�&V;�8וqD����朡�\�Tq�1�����&g�kd��݉�
���H�(�L� f���*kK�Gڿ���DE��r׏;��p���SI�gi�$�x.�5ρ�c2O]��5�Y�;���7m'qg�(b���i���׳X��"��[��Qv&i�y��}jUIP��~��(���
����Q��0̛����� �`���s�8>��R�����6���s�����AoF��>��A��ap�_t:݋
0��d��$^�+Nw�l���TqR@�'��=�輁&#�Vx�n��q��3ئ�xc��r]�C�ʡ�k�WZ@�Jޠ�Wr��� ���y�W?yɿ���g�zk[8*�3D�uHR�]]�6M�'W@銂ղ�Z	X��R���8�V� S�Q'����G���'4�����ͷ�OA�����)���Ry�q��Pњ�Nǟ�ES���Ť��������J��|�Ɏ��*j��CN�����a�%u��*ߥ���_NX���e��4�j�4�v_�?jJ�.1{Y�0�5������w;��$���e��(�V7�/>jEnM��3���e�7�G�� ] �L4h��r����{�%Xb�A��dk�6��#�u<-2A%I�� ������/#~�O�]� r���׏ڋ�.�=��h�~��旍�_�3�;��(����;�����H�EԈh˼3��M��$
FO:ʹ�붃�}V�\�)��XZ(��ĘG�F��#'�4��%��/"NO�0�d��Z^`;x���$�Ë�ϐ�G(�tQI�@*<�{ ��!��"@�b��� ��4��G S������~��iD�eR�v[��?p2�;��h�PG*�K��?���}�	GhB*Hq�_>Td�D/)�C��]=2��id\��
q��nV�5��.�v2ĉ��X����.�~^݌^��z���ƉKPL���f�ދ��S�kt ��0ݥ��+���z�Ӡ��Ӵ�I�RJ��{tw�Oj��Ѹ!n)��]T��/����I+�w�驶�&ګA��\h�>�;������1���clZm��4i2��=�h�ymF��t���м	���+��q��ީ-s�i�5B/�v)b=��u�~t=m���'�\s���q���/��M|�kS����̆[4ґ��ֆ�_�3�f��lR=���t���ix�|NB�}�&��π:�Vf��C��S]g��W�#�ڶ�{ּ8�[�AҮ���i����D2n���Ei���>�8J9#�[�����JRЕ�Ѝ���lm��o[�K���Mv�]�0Pp���A�Y�gɰ�1� $�*��U�� p�ag_Ԕ���Dk̃ףY���x��2a��/��<�ҟ��(t稘��L:������vҕ����tR��'<��`$������)���z�l�1��݋������JҨ���mU��g��uS+v�RR��ڽq6R*s�X�n>z9�뵻/fon-����~.�_�����ٵͷ�6d�<"0QMnZ�')��2 ��]���=�%�'2{h}�GE���]��̖N�#���vl��������T�[SNҳ%�Ćy�T�����0�֯˽_b R$�:Y}u�L�	�:`��D�%���N�n�Sݝ�&u��)iIt�����g���ӝ�)��-����ל��1�H�?t~�^�����bvY;Ѧ�@L�6�o\)1R��m�6V��l��F�CH�JǍ���܀��MBr�~���Uú96ս6Դ��d�RU����T��������7<��~qѳT�#�ƳD��^Ձ��T��Uo5%)�D���8�fU�Θ���ƐNW.��{.=A���"��[#��w��0�Z]3_;�#&ޞ�s�"@��-�D�&�����!,'i�:��]��⏐��vߦ����=�� ��h����=�	��y[�H?P�����a*��#����ĕ�0nH��i�����E9AE�.3�bx����4�z��V�[T=z�XK.0��4���ٿz���HeIT�Z��b]D����+&%h�\�_��vm��e3+b�*>�Q(�~���K}�n1�Ќ�ԊJc�՘�!����₁͡x�:O&R���<����me�� �ĤN����'��2e�{M�+Xuؽ,G�).w^d_ilT��
��މ��ѷ�|�&4n��~"4˛���5�=̼�<F���w��!��w�<--��X ��۳h@4X��
�qC���#>�+�F�/��L�A�$�y�ьZ�}t��}��O~'߻��Ne|�I���A��1a<����!zɜix�k�5����|�B\�T��I
���k:s9"g�U;s���C�7���Έ��4~5-�f�ß<P�ߒ )L3�S�����w��[E0�5������)8ؿ��3��/ �z&�'��8<�� +*��c��k��qj!���o�8����y�9)x��i��M
�Ϫ���R`_d�}�v�#�YYד
 ���@+�����|Q�,�/���YY�2o�[>=dmI��E��P���oMqe�Ndl�k�H��4��t�I�{���t�F	_�������^ӕs˦���`�#��Q�����LV�A�`����4׏bR ��H"���%�(k%�?ƫzg���	y�\Ӝ��c�(�m��P��T:�6	���g���m�a�������r����<ɛ�\���
A�.��n����5�P��t�`<]��a_�k�QQ��Dh���;F>�g���bX�m�	#���=f]UW��o�	�sj?��j�;/K`s�h��O�����r	u���*�Y-rm���P1͚�ċͿ��MΤh��5�7�Š�9�-�E.�����T�Ot�A����TaH�!m1�^?��>/UMk�b'���W���KP���)�$�U���|��,��~Ġ����]���ty�	g{D$"I�ad'Q:��J)*��-=F�k�k�E�R䴹�3u���|�y���1�����G.��9D���[�6J["H�ǒ[��먻��AG����}yA�ЫW�g0��b� �ƖF]к.�n۾s-�LŚ�W ����~�ۅ�\�,��a(�t\�du��w7�O@Sl�zAbȷEʯ�Ȑ'3ȟR=涄�T�H#S�f^h��R΋��t�� ��ēM�l�,��9U#+H�:Gt�k�SIB$� kh��Jv���S8�K�vu�gǢ�Խ������[�w*F�F�"2�?�O��k�qҠ����1+L����=�<C��>�+�F}��(��h9E�-p����&�9�+���_���Z0� 5p�t_�B#�M��c��¨8�t �U�@�� ��,���
�۸;ML�E�[78ܗ���?|��l�X�+�ü�T��A"�L<��G�?��9����G���K���QƑ��O�eO�Rek\6k�~�&?�@h�;tG5�Qc2`ŀ��4+���]��uS��,��;?�W��(����N�"Q���֨\����Ԯ�C��)���̞M�g� ���_r�g����o���~�)��aÍ�AlQ\����yw��	�u���Me32
���}����{���I��09��4\SX�&��pOe���E�>`����nJPXZ;��|��k}��@+��x����so%��������8�vU��D��-\�hZ�n�w�	:W���������)6��*U ���)5&X ����������c�g�����yu��}Zʹ}zX��Ҹ5<Z���wGeb�7�D	u֨�eHp�^ƀ���J\���?��[��C[[��$�܎"������auP��G��#t�JCtQ.�z��%�^�1�>����� m�=�J��AEz��՝�]������R!�]�2?F�>
�?z��t7�|���f�)p3�-�,s���l���C����Y�չ�?(lsZv%��=��#�]�����S\�lY#�U(�,^\�/�s��h����'K��]�}ڟa������p=�2il���q�fVk��W��/+^|��� Pg3Dŧ���>Bb��QƗ��b�!^Y���O�FH�!G3yΕ��m�k��%5��܊�,\pc݅m���l�*j�k�j�效_QM��c}/u�ZV"��n�%�+��Y#*�v\[.���]i���B�,����'�uΜ�W`
\�i#����&���B-��.D�kY�gc��X�NII����gH� #x�j�Z����LRps��#��Z���+���e�`�(�o�!L��K���!���~�\�
����+uӰ��J�6�3�9{�]W5?��3���y�hb?��}4��;�3��F3� I�p�����9���s�}���\�"�ޞ��r��]�~ h{��}�^k�L&�ZT�[`�F5�+P��eJq	H�z�Cm�f�R�����Q�t���2�Й�4�۠ӗNs�]�{�2<�����PFl[U�)g9r�tgW���|ۣ��~�ȗ���~�sX`�Y�,/�1S�4��W��o�b����q�ҽ^8̭'A@�gN���X��榠1�%B7nC�{)i�K�1�#^XL�x�!ڗJ��~!�~V���{���;�	�*c�����C��`P<Qdk;~�E|��V_C_4
���a�h۬�W�7��ͪqD�����ց�GܯP�O���?49�e)dFC%��_���MN?�C2�n�a�X9]S�����sq�i�z�%;K ^%.l�p�h%�1��_�;p�15�'�ez���f���Ϲp��$;e����0��C���&.�>R�s	����{��&�$n���v9��8x���ȧ���ؔK��1��r���vH�{@��o>F��d��r�Ơ>���u�����c|����LႪ>m��qG"���Y6�O��ҪM)�ha��
*���v�*/# +�W슼0蠴�-�Ć�ѯ���p���3��;��5���4�d��\�O`d���ΰv1�fm�J~M�͢�l�< ��� �t#��?��-�V�a�i0��ZH� ��L+��~\��P��L��c�P���x�=֤����� ��~䙬�YLI��	{�����}��~���3Ͱ���/��| t������^�O��AUL�@F^��N�0)^�2[��O���ZA��5�u�[�	����D�lB0/8c|n��k�@�ik�L�Oz�����E���40�L^��?����y��E�X`�~���<���e$Ô�eb_�X�K�}T�|��;K��.ј�=�t���#&���Z͚�'"��-�EG"$U���aZ����NT�'����_WE���}�|�O�_[tK� �#HA%�ç�\�5|b����6�)��z�A��;<��륍6g��u�#�n�C80}�[.�={A07~ ���x��TS�Q�hű�0�͇j�*��x�����r���4�F��|l�v��z��ސ� �;0���E�¿����u����5m<�`����z�zP�8�l�ŝ���-G�ĖUK-G��[i]dJ�Q~����� �L��H.S�VV�(�a�ֈ�o�5�Cv��܈^R��;��e��ϰ(��r�j��PPT��翃����!�|�	+�*#
J� ~ah��I��T�d���=s݂���h����:H��Vf��*4L��U�}\%kax�x��|��&�3rg��B�	8�W��%����Q� 2�:�|�9G��s,������(���V�b�7�m���/X������*?�"oR�s� ��l����c�׎��kRsL|�ڷFW��ƶ�f�	������vj�L"���d��Ӭ7)��Ƛ����vay�x�4_y�n��jS���8��h���hu_�����.Ά����AC4���D���M��tE�i�����#��`ض?�zm#�Q�oC�n�5�>��C`��tƟ�c�Buɘ��e5����[��6����S^�?rhU޻E��[�e�-ݰ{m�T��.֥����!1E���[.��c��jU�(tݚ�;��
w$��)��/I�	^7$^���#�����c6u57��j�Jq���8B8iz^f,��K2���`�lS�� ��Wא�0���}��u`g�W��2��{�ʊ��H�ą��9(E1/�L�ﵟ�@��S�W������On�1/��*�!�r��%�FF�����)?��JC�zF��V�	M����V���'�����䨒c(U���A��S��o�-�Y� ��oi8��xX5i���<������fut1����jV{e9�\J�bb��J<�ڭE:�H`����AH}��A%�91���
`��f_�V�ImOU,����cqAפ���ɳ����[s�լ~���Fg/<��y\�����4�%ז�SI��?���T�Ч9�e�>bF��L�d���1h�����p"E�]��@��Y�Vf�f[��8	ā+��L�R]<��t���{���v��ȍ����DK~���Vo<�
ݬ7O�I�A�"�ڦb�3� B�%j������ń�+��$�m�Sq���[�`'��iӗ��fA	�_��R-��]x.�.-���q��B�Pn�~�Ӽ�eP!���&:�q��<][���B���F��:i�����6���^�^�����v��/'���w�.���@�􃺜*��蒚r5h
`��(K�3Nl��Մ6O�=��ߏ��3Aԃ�J@YP	^�[i�ݒ
'��G��9Tϙ"��oV��c$6����݁˳�4���p8���2�L�с:Y��C�'�7jC�P�X����DN�h`���˻bN�_ޗ�Eh.#lw���)�R!�&GKp)��l��WP.t�ZFk�MR�Sx ~_��#V���r����<��{�տ��:/�t?]w��(|�v�
l+�V�ce��U[")!h�"��{>�C(��˗���vuX�2�����	i�Я�2LbB� 8FZ���`��~z���]HjQB�A*�h��Z�������ؗb���]��ۆ��R�����ߺy(���fC��`���)��?�W��:�t�&Hd���G�=��W��~��RZ�0n�O����Q���v�e��|�-~j_����'!v�A\��y��J�e�
����*kN0)��Q����e2�T�(��͎v�#�t�����Y��QD��=�P"�đ���� ��B8d��T��ӆ�¬<{���1��v]}>��C�^`���nr 9�?񻞾��u��Jxe��wSs�s�Wf�ƏW�T���y�񇸜���+:�fg��) ćb�=�	��C��@��/[�������i Z"J�r��f��5�s٤�?�������M������yv"��<X㜾9�4�#�sC:Ta���`7^,Z�:���ZF���ܿ~�=���'��)~K������4˧x/c��h�����-ܖ#�g��j�M�F��sn�;T�%��1�|yL���p.�ʣ���~���Q���q�`��(�aQ(+z1\=�
��f�"���([�Ϩ�p����}9�[Ff�B��뎰�m�j��0�X��4��V+�h*Ä�����Kl,ƸK�<����&��>�����,�3�{!���#���5T}iD-^�*^�UK������6*���G��bn�[Ku{M�Ut	������y=��칳v�Z�X��Pb�����Ele��ff�@?������7�Y+�Nq����\���%3��h��e��[�0O�����T���6~}q
@5���E�λ�8Z.sg9���@W��&���&Ѻ�N? A�>0~V�3Zb��tK섬1��*�'����JAG�)���,qI���z �Ym�� ��ȯ5�}7����ͷ��a�,�8�y�s�H�F�3pU�`�:_�E���mɌs��7Q��@���;tic?2��GœRug��"������A�^��� �������
�Hq���r��o=��ZaH�e��Z@�F">S{E��M���B\{�2=}�{�j�2���MI��O�:6���A��<�၍,�5�������wA3�P��/h�W���;���Tz:�ψ�.r����S`1�*-��!�HS�H�x��$j,JN��B�`kr��u]iP<�3�A��/��t��vήP�n;\�z�[<���5��\Z�!��t��4�4�;�,�S�^�fzuQ 3����Я��MUD�v����Y��B��U9��C�ʹ��+��]�?W:[��:+_+��(�B�љ��2�F�Y���N�4�Q��f��L�{�<���3�e���HJ=۸�p�d^B�K&�y3�5�u{����M.�=�_�+�8��?��I�GG$�5�������][34X,�E��`G��6��U���T|����%_s�ګ(�0�֍ CoQ*DS��5A�܉��Bj&���f{������X e����+*�@�O�^p74FJ��_�����l��p�u׹������s��8wz�#��Z�<^
��^�9*I=��0w�x��d����%�t (���a�P���Y��������Y�<L�����sSO�3��*!�DXh錄���4S�YĪ$�&�?��0pi�{�����ږ�����j��|0l�g&�W&� B�y������p��A5�Ln��F�!�ٱ1k�w���e�\
�c����6-�e�*�GlLd�-|.��O��ݏ[a'�_M�΄xؕ%Jџq�j���:P?�`��.�O��L����x�%�r��"�q�7"�F�C���&~�P$V_�^^�3{0���{��"�X�C�뙵T�Z����	=޻ժJ���B�'�h6`i�&)}�7'����
��)���p�$�$ۡ���i�"��Q�k�ھ�l:���,�%X��Y��H�6�r�6KR)�+�
w������-�K�j�\ꈵ
��F� �eKfԙ�ڥ3�hFIY1���t�q�Jr}VB�	5�����8�9~�w�:����F;x� A�o��A4R@�^τbö`3x��h|���w2(�a8�ՙ4��G�:�g�}�W��5�u{[p��k�ܰ=����A�ש{��䅾Y��*��0���!���Dz/�ڛ�;v�<U�~���g��8��gBG���Y������o�S�D�\P���&4#̘�o�b�v���j�뮛9]�p-��`Ea�qB����7�� \�4�YPX�+|;��{���ƻ���m�#�����L$_������:C�wJN�ֲ�x�|��Z*Ғ(+��:����s���ƣ�XP�bj[�\�׉����A���ᯧ��**�&��:G�4����c�'��������O�;(Ezљ����\�/L<Ϧt��n��O�%�2Mx���V, E���>D�^��'���H�Jrn�\'Q��t��\�d�L�O{z����Ti��?��1��,��]���s+~Q�;��xDA�+:oӞIR(���^����h�ψ��Dp|��?c5$JX}���d9�э���(��f����]	���]��X߳��i�dy��t�Z���벆8�ۄm�,*�b���M�K��W�׫��*��![cʄ:;h��6�1U;@��s��a��a��n����|��P���Њ�̃��KӢp���;¸�Y��H"��npE|�s�����O��^����z��r��� �D}���w�&�(A��F��fF�ƐW"�V�k�k�@��\C��Ɂ��]Mf>�b������J�4�T}�2�FD�H�0.=0v2�O���[g�H������T(y6`[b��EEU]�\-�$(>:?m:+�!��];2�a��f&X��CI�,�Xӷ�A�ux���;�Q)kؠ�x-y��0����词fJb�f���A;��|��:��·OZĺ�ݠX�|�� �@�s��Q����C���]=�t��b�����c�H)9�����-1H�& R��|maS\�k~/4��?e_��2c7���u���o[�?���_ڀ��
$Sxi~)�ڹZ� Vլc��n�n�`�D,$�ڛ\a���JMF��.
scmb������n�¾�,,����XP}h��3�T��QY��a��O��פe�\,.@��K`9vѼ�0H�т��N?"���bjO&>����pG��n���ZX��aM�3��H����h�|u�֔7;���h�nK|��C�\��y�����Q�p'۷�Aj�>�F!�P���k�y���UD�ez������vUDjb{������:�Wi�nF�����T�F���K�6����,Ɋ��s�aZ�*3_��>C���` ���m�m��捱��?fd�A�(�uy��|���������

��`s�g������[	,��$^�;2?<|b|��.�푤\'�?&�c��8.�Z��x�m���*�z��=��Va���_2�|�2���1AU�ehr�E���4��:�����D�L>�
۸�}7��v�a�S_�V�V"��/�O\��/	}������j�*ʗa2
V���]h�|j��h�AAdG� )�n�]T���5�~0X-�A-e$�Tƈ�d����͝K��-T�ЁE9J� �]�$MG���)T�.��(��(����N�	¹�h^�����zHUBžQ����M9�̷oM���ϥs�d���,/��py�"$o�ׅ:�}��.[:����;�CD���ΫR�	W�λK�rtP�w�Ac+/��+kZ�y���DOX:��"Uinչ����Ko8i���L�I�lg@M�LC��fe?^�Ǥ@P�L�� f݈�3bm����W� F�b�'��GU�cs-˂T�F������/�����l}�8��ӱ��Ֆ>�z�ѥ14��K!�s��t+��>�@Vؿ�V`:#jk���! Db/^��(Ô��{-�W���{�ͨ���#xd	rwH��π��xm�.������im���`���9y�Ë���Pt\�?۲�"��UwƸx|����8�����=D�n ���\|�iǕ�n�[�dU���*��+��o�����9�{�8�I5��jȈ;����-�i�
3ǎ}&O�NkW����A�$7�0/�da��M��~�X���ڼ7P�8u�I��ÿ.r?8��W�a'W��E�p@hZ�����Z�uo?R, PU���.E���в!�A.��W�G���U���?�X�zΦ��c���SV�B�cK����Z�9�����%�}T�c�� GN!�|p�'�c�:������J&�`�C�HϜ�
�z�T�i~e���o�F��]Z�_���qs}��&_-d��U���ޠ�H#�[O=���^4s��E�7C�%Q]�]��qZ)��I5��}v3
�|��:�wX�M`�5�CkOf�O,�������z�H�B��v�q@��(%vL���~ᶔ���N�Y��?��6>	D����}�@�X�S�_���^$���5�7�'��B�	F͵�X:p���� ��4�*@����e!N2�䷣�;&����SdE���mܯ���)�4�J�h���c�b��:u2��U/�˷m��e%o����-�c�o> 1��zR����m��������V�U�0�������0�M��"���*��7����
�
D�k٣r��e*�e)(�f)e�|��8B��H��`A��"��&y,T�1��'�u��pe�h��)n��J�/V��C�pa�8V��ɧQ,ʎlk0��r<��Z���e�S�s�Z��b�A>��r�R՗�&?����bq�X�j7��v���WK�J0s%tD
22G&�� X�K>�|P:�"�鼺.#��厴�����o$���N`�d�ݏAato���"/B�s�n\}?g��Rǡ����PCa����x�~��٭���QL�	K��!Ii�nov�z"���͸qm��������]b'R�豀�%x��XR�x����*���D������>�sFh���)�}����u�/<ᬬ.?�%�a�zS��ds�;w��N��a��oh�]��`�xZ���e��y�Sf9d�F9J���k%꠮�O�>��������(6��Ov��e��TW�=��N�Z����ֹt���m�BXН�K��1/VA�����ׇ��O&��j�	�����7n��&�k��q_K�
�n7�G���ΰ�l݄,3
���vb�[d�.|�#39��J��X;1�0��� * �-Z�B�s�r�{���Z��~��Tf�\cJ�daa��H�.��*��)�E����bM�&��c8�"��w����V��tU�}��CH�=*P_g�шj��ל�>C��C�lN.e�Hc �����]��R���UpҒ�=���OY�_�����%d(K�}[�~���	8���T���5��9fe>O���y�E4��*��`�β��Ǹ	�5Oj�_�M�z��!Ǹ;o�0x��F�|8����ٗ�������ǫ�ơ�R�#ǲ�Y���(�,���^L��!�AT4��Y�ޛ{�o
'5�U
��Ȼ_C������5�"����}W��.8��c�N���ލ2��k�jk�a�����eSp:t�-���o����d�ѓ(��\�0 s�6�|�ɔ؉��Jw��❶��KDq�sM����cFk�-��4*�� �����T�B���%�3Ti{���G�*]V�p#��_hE�0^i�ew���1^��d�}_N��D�#���t}�{���O����{�#7i��`�n<�˨��i��d@׀�+C��X�\~�{���6��!��X��ZL�dBL��E|:��Q_R}��V�����3�[΄�[���l���	�ˉ{<��q�#�g+�UC��ZVY�	�g�d��3��(��eˁV�,#'�I��$D�����@Bg���f�H�1D���ߒ�1[�j�͇�0�3�e��8	��m�_?i48����w�Ŗ ����&����o|M�ZT���\�M�})3&�����
����+(L=ar�M�v)U��}���<��L��߷��N�y�,�a�l�����Gl�I���`$�$��h����6/R��/}��~�QX3��"��	�G[�'�#=z%���'j��XA�%+߻Fd�C|o�૲����S{��"�U��Tk���S{>�o�/<���3,���=Z��r#nS��F�v�#QQ�f>�f�kO
U%�z	��&�l�'e8l��������
a�\*������#x<���8cz�_}Ivv�|�n�� ��av3�wD�(���H=I���QmҲ@@Mz��8ki�0.g�pMGi!���}1K��Ү�`�n�6;��XH}���w�X����T8#�γ���bܧ�H�D�p	��ڂ�^�K$|�K���5)"�1-��Y��TW�� ��Ru�=�9 p�s�3�4=�*k�2���@e$I�X�)���+���4K8V��<&Ҧؕ�wH2v\�iO���h�U��iϧ<PΥ:y	X.�o��;b!��!dP��ʄxM>�=i~�H���Y��U��?u&��Lb�\C*�{�P��(aԆ*���|�`��?����mR��U�a��z5�	�H̠R��/]9�i��'��4;��5�>S6����p@b��#��x�b�ܺ��d-Y���<m��	�L�x���m+k�P<�gj�	��w�����:��M+e�,�����kx����8=4:"MQ!�ʐ: �7�)L�qn93kg*~.~A��H/����Bm�igèlm*�-f�>���&�2��R���PP��O�׆fc�H3+h��F�Ae �[�����P�E����7d!�(���^ k�7���Ļ�vb0���D�.���R$�}��[	���,ڒEf��`�ᬽ}�/T��}����3�ie6�R�']�p�T��ku�# L�/�Ԙ�I�X��#mU�H�}fdWޫ�}�-��
�,��%yɿt
�B��J
du2��@��Y<mg r���p�"o?�+3���K@k�ؙ��В�sC.;ά[��=�C�2&w��b�g1/4S.�����k?8������J~��k���m�$�'�f2n�vBq%�X�c'�&���I��;�`��!r˙~� �
?<���>�>��j�.~V������"���>�Q�,�I)L-?�l�
u9*���agb��	��`X!�r�!}�Z��"!"�]�y�@/�.#@ Ej�Zmv^�%o�#�W��?=��ae�-/V���ޑ� ']rm�;�&�5�@�УTͳ�Q��c`�oT���չ�,0 ����Z��g���Z$�Dq cB�ֳ�-��(����YS/��"@zTI���7-�ӿٔ_{��^-�gCH&V>e�����񨯽���ҧ�U�q�r�M�?�5��b�iJ��5t}���i볏�Η�gl.������Vd�p�q#n�|��n���$���%q;�9���-=��gu�`���{`,�-\�?��'Ն^�C����Q�S<S��kd5���I��\�FU���rL�9/ZRO/
�oЭ��)�Y�C"�+��4�E��?C�Lcn��0c��F�I����K�A���|���w�\�k��HvV<Ҙ�_ӵ��#Y!��l���ā05jK>�k:(��*�7��M��a�>`���&��������	�sZ��
&QFn����e��۷>$yL�a�;���VGB(�|�^���@e<�>�]4��R^RN\o�O�q�'�[�K�B��eG{b9�Q[�l�7]��L- )�z���m�蜏��Ut�ˎ����fL��+�"B�'~b5p�'>�tĚy��������(sY~"� Dc1�Q���'�B��	q$:����ڜz���ؔ�ཎ�Ձ���q����N
!��9�3?��-Q\�=���}:��R���Rk3��%}tE-����j�C���|����������%u�p�ɋ��c׹�S�N
0/Q�y�Tf���;Q[�`�R�-�
eG�n�	� ���,m;�[s�\Ѵ�4�"!_���3u|�*�/:9��pZ�~@o@AP.,�$M��8�p>��bH��b�h����#�[�({!��28<7���k��MZ��_������+d;
�	��%�Ty�~13��,&:Om�&"�z&�Q<���	�W� J�P_�����-���p<I��&�d<���)��q�+s���꺋���q!2PJ�t���e��,�E��cBWԢ<&� 帑vU����E��]\���~="��4L�V�"Ny=Jv5& k�1�f��9cΥB���y�¯U@���9�,���9�Oa�x %A��b���;e	�|���9Pſ��ۚ���]��;�Efk+(H-p��%z�Ɋ	�sE�8$��B�����\[Q7Ş������Y�+��u���?��J�a�.��
��/@� �YƓ�[���ӵ�)�d��%9���o
�����`S97��rA�s���9����	�����~�'\\�al�-��\k�����W��t���u��W��9Tj�&p߮<�0���=x�⏦��T��3!���i2��(B����q�����}T�5��f�O�4Kc%�aF贆"r��y��:���E�vY��'Ƭ�Z��D��[�$��4G�re�;Ni�zm���y��n�k���������c�%�ۘ�qt��8�Y�7K��Y-KӉ΅Pn{ئg@:'���*Շ�C�(�QX"˽�/䨢��͖��+"T��-;�� 3i�s)���w�z ���^�|5 W�r�`K[_%{�b���vP�A��>-�g�aG�߅[�}��)�g?&�U��&�V�F�JbQ?��c��i`x��,����΅MLoƞ^ШS�&m��� ��Z�y4�_�2�1c��,[oaa����Gx�(z�,\�,=j ��J$��$��)���/oӶ���Y�/J�+���������]M��v+x}�nw҆���N�Q��$�i˰�@�8+f�1�d��
y�{���t>X��SM�f�@ �^�#v`�UH�:fx���8<�F{CO��|P��=W�����c� ���`ds9@HzӠ�:ieә���[�|I/�� ��XN�[\�$��W���8R&�S��������̹
���X�B�H3"���Ӎ�2��]�B���si~��}񪮦������r�Sũ���K��}���$3����T����YAΆd�(F� `i�|n�"��F���vR�{m�rqb֫�|c@5d+m�%�Q��q]�!߂b�&��?��Mݼ	���Ė�J�(ʑ�#���0+�C�FNgF�=尢�A��+@tgp`u��
5$m1��N��]��<������r���٦>/o��|� -&�	����]a�?�U���{����.�b����]�ץa ��K�y�b02P�A����\���B]4��_~ �?��q#�R��RڝZ��mrϺ>g�����ɳ�}��l��R����.+:d{;�J  h������� *�x�H�H�
7s��$rL"��t免ky-n]��iIQFc�+��&��Ƙ�bPD��ˢK�>e�ܴ�@&�-����`��!��0
�����'�$m/Ҧ��D�b?v���;���4�@�*G�߄��*�����J�IC\����.���\"*���R����{cƙ�M�����Iί�.����p/�eG��C��aq�9��F��r��s3�>���s���ݻ�a�Z��_�� E�;6�)�P��<�]!;�|� C�P-�Hv��ќ%.��0O��;���cf'ԧ���=V�Z�.�)n[45�rW�X4���]G�ɧ��Q�ׂ�_"�f<���qJ���O�~�!᫭�:L��Y����_(�~1�Y�vV�_�SI����	��7�>٥u�y�>���r��)ߢ��
Ё\�O�zݞf�;�7��y��:�
^*~�<=d��^c�.��-Y�4���kQ�'��0�. +?��]���t���Hڋiؤ�7~�B�i�n$�SP�y$�0�)_���Չ�O���u)�D��;dF!��g_�T�kZW��@"��s���Lz�=�Ƴ;�-e�d��t羼?�e���V��1�����BYZ�d���8�p��r���D��hx��襎�
A(6����-V���L���k�#���#,�}[�	�r]�tÎ�e��J%R�ӴjnTF�ݞ]��E�~�[��䘒�w�1UO�͇R��#
�M7�tZ�2�o��Xf��8/�h(����a2󲷷�)���$#�o`�(-�v�m^�/����
+��D�@r��ڪE�;x�l^Bj2b��i�yzJ*3'�M�����%����^�C�h��И����q*JTJ�}Ɏ�~��9���:�U���7��&�� �''~Ef�2�vn�p��-cP@�!M�FyG~X�m���u_%��DNH�C�K���\(�@��R4e��l���X�XjXڧ@w�dI�������ј�ja6XX� rV���pETqhn��Q��UTMX�!��rJ2=�)o��x�a�LA� Y����bi�a���}9���;��L�_�mN����>ȥ!���\C�]!�j`����77�	�����f�Bf�ٺ��
�;h��ē�2pMǙ�E������Wjn�0]Dܡ��"�=Ϙ_U*�C0f+>�ɤ�ٽ16�}�� ΐ���Q���\�}z�*���TKCs����b:�#�鉜ܥ��;�l�j��+!v�����Ic=��O-�4z�NX�o}�eer��)�G��C����l%���[������a�(5���i$����i�w��|8Z��f�pE�0G�X��	��C��2��@�<d~��[G�]�ĩ`g��,ˣ*,�f/f%2;_�$ʫل�  �W����j~(�������Ŭ`�Z��I�@����R���I�m�WH��d��2���iE
qJ�N�R��ːI�y��ipN�hy�0��K�����i��O��b�oH����Vu�J�Ѥ
�\�.��7U~�7�)��Zc0��]tk|�?�`��-�&m���Ηk�=�1҅��'����ˬ@�M(�¯��߉G�-
��e���^G8ܡ`߃���)�{��94�O��h�� *�֔���K��=�A�T�_�3�	i��J�e��ʐ�!lh�MlJm�����Lefj���&�}@�|����W�9��ܱV�v��M�pWps�Q�貮V	F9����,�(n��L��C8��S$���d.�k�)[�C��Bú�Vmx����"�Q
�D/��K���M�I|A�f�1)�2�N�T��C�F�7��d�_'��t���B�?<� )���֩g�:�i�8�I�!�mm��p�Ԕ܂�����D�30�9�-^����L��խ��1v�͸-��P�̂c0x����C��[훌�y X���aFDEח�al
uʶvSo���ڭ����ճS�}xR��<�%��x���s�69��e�'�����C �ޛ�d@:{�K�+�Ӯ�f��>q����?�:��wzR�m$�����9���J�tK4�S�n�!1Y+��	okx���@rGl/inF�lY��<ߟ}���i[���|�+��B���䃜 яA��+��C�����:��I͜o��L�D�."CZn�_r�KR�<��e��'��8�����h�p�L"�T���v�?��t��&[<�cp�刡N I��s�g.�K����9y���̷�F�#��ş|�W���1(.�qP��J3K�a���V��C(Q:&����o�|��ͷω����u������ee�
��/�~$֩p��I��c>n�d�ڳJ��`ܲI����VQ�� O�H��|���pI%r81�8�i_��ׯ���S�B��j�ڟz�zɊ�r�p$J������z��6��F���a�fA�	�N��6R `Y$��Q?K���/!�3F��jG�؍�`9
��2(��� r���*�r�G�b��ش* ��1�x���A�ӭ���1O��eZPd� �������U(�D	���Y�1fmt�VP��|��;�V�87p��;]?��+"�Zv1�����v�%:;���W�Pv���J\��������1�U����ꣃ;��@���0��jATM�1���{g�liP���J�u�:'#S�Ǡ�K�uWv~��8 ����HP|f=�щ.A>��İ��A���ԂÏ�$�)!���6�|�#ό���h$<�JJT�XĶ���@/N���.wev��$����*�	�@J&�at�6�L�RS!""���,��p�_���L��>&��Mlܮ�� �ўr`o�b��L���):O�S'�9�gսȢ�"ag�h~���'z�s��sU�G0�X�e-�l��#逭i�,l9W��F���v%��6T(UڅA�TP��?v��M�x��'KD�J�,0�	 9�.�m���'٠�M$���i9�=�J����L&v�@H�������@s?6�!�[g~�W��)�Iۮi�7��~�6��S6W�<R�e�o��q�uN?M[��������Q�C劈;5�����J�5� J�E���������0H�����$��� ���Β>���0�yÁy��(�2=��Jc�)@�Pzx��0ʖ��|�f�v4��4"����0TEs*i�;X����n��3�a�2�`�g��dh���?��W�ħ�2 ,���7y�b�5D�H�K+3�'w��Δw�����#�5�\�k�k�k�,��գ�����***���Z���m�Ct���OEE��q��kB(e!1�~�j�,�"�����O�������}_D!3���VO��A"xa��N�w#�Ǿ����h��S%�|F��Z�� �	�,����߾���h��q:h���0��
x�9��~�\���he)L֠�89I52꽳�	j�7|8 ��H����'�G��by��ЖW�<���@��f4-�e�ۅp�Y�B
���a'q�H�0���>�P.�O�j?�l+���<�m�2K���7A��5�=����4�D�G��d��r���s�R��/u�qw�?ؐ���s�����T�8�C�q�tm���,G�'"��w�����w�>l�A-́�=L����3�������}Jm�B�"���������T��������tN�`D�oP����҅��{�Ga���cG��	#"G:\#�$<��E2�~��0����=h�Q;t�Ê&�A���#�~��W���z�]�2זMb���n�l����1��خ��$c�Q��"4l��;\h����2t��pu9f!D~ŀm�٢��f�kq
�oMܛR�l��3v8\��!������_���r%�0�l�&Wm��ua�_z3-�,�6%���D4�����9#��3}�<fȔ�D;�_���JO�loF[�@�^���憲�'�H���~P����P�O�?��	����k-����#�O'8��L���.��M�#�у���S�b�C�t/b��"o�(����-�K�1�:�U:98Y�;��w��&*�C��Ϸ���p8����MT���Ul����xy��� |�W�G�d���%]3?7�w���?�b�k?�Tg��-�2iҹ����E(��=��o��u��4̆s��¹�����i/�^���#�k����b^;U�C��Pa����t�U(q��Us���%X�}T�����zhm��|\�ҡ�'�Tz��v���)�+L�ӕ$̭c! AQ�(�rI�� �mɉNc�����3�b����Р�E���T_�-2:܅!L��(p�8I�M�?�9\��;7Z��+�&��颺���y*�6�/�&�:t����#�Ɛ�����T�2&��RgǨhEQ��ު�S��=��I|S<�@���X�x�^_����n鑯�	�RB�������R�W��h� ~�K�P�Q��C������P�T>o����!�ꕮl����������T����>��2�l�ڋs�:"j^s%X�9D��C�W� ���/�$c	�����A�hTO��N��^����n�G^�DO �\53��z�:��g�/�u)9Ə�N!�X���ұ&/(��NV7Nm1 �XT���;C��M@�]/8�L�t
H�NM�w�Xj%b���]ϙ�,���\X���x:���:����ˎ�bd\��>��oP�A�a���-hlV���0�M�I�c��Xj*�B���Pyy�җ�\��}!{�u��	t�\H��n���>ā��ߦmL���ɘ\��P[	�k�[7�ھ�+]��^��'�D��q�Zq����b|��R�fk�jr�9q?��gHf����H�zѵA�L;��nwCFW��ǝ&��j��a�wMӡyEf8A[��k^@ʦ2<��i3�ݞ�f?A[��FD>��Y$�(X������.l*v�m�$&G�I�9�s"Q~�JѼ��fί}��R�3ߧ|�j�ǖd�!���#R�_&e��Y��;��l�x�����%�3c�ʃhwf�C��O�$4e��[{�cr�SO'd�+d��Tn'�,�Gr�E��p 1Xq���~��]����"p���sΠ�c�h�wW*N/��2.q8�d0�I��[U��jfcu��7�T�Ư���.�j�v���-T�X$5sUͬfs�O��.`�������o�=	ԧ��`W�R�/�N5���<a#U�	��?'��zK�Nه�5{���s~'�?rS0�?*e}��m7n��r�	���{�?�����7��S|��Ԓ�:\AŶ�P�9��|MX��M\^������2�}��Pq��[+5|˼���
����l�KEc����^�ܰ��G����#�NPWƼy�v���ּRQ|Ql��!4�f��iȓ��AB��<9<�1����=�p� z��O����1�� )԰P���7�2����p$��6�r����){�8$ߐV��W������8Q�@�� ­��$#]{����H��\b��s��$A�\�*�锱_�#5���Du�<@^z�ƕG ���3K&�J����b�G�-�� A&'�nƫk�� ���8ŀ���L�L$~3�����nh����eM�6��?v����Q�ב*pfDC������Q"�5�{4���4��`|[e�d��cO$`ǡ��yq�ȍ�2�>�'T��i4��A�`�:�t�p$4�N�{���y@�O0d�Eqd�xŎ���s��oz�+���	񹈆�D�/�)��04���M��͖h�O���76;p���C�éM���0}�B�r|-=*���&?4K�M��T'�}ܝ��"�&��%)��M�q�W�w��UP�8�K�nb�F`f��Gc�����ƽWdqn���b֮����{bI5ոjai�z���c$%��$+B6��2�e�T��!R'!�D�>R��6zZIRƟ�W�5q�'��/����Uf��΂��`4$���LU`qP5��집�FV�J����k6%B��Y\�,V7V��-�����.{�H�)a�2��}��>g�ԡ���*d�jw4�Au
�l�o�m$���(�w6�`"(��Ĥ�ǆ��)�4�t<3=������3%Z񌵋�V�%�t9�@)�u�4�at�F���<����7��T���5�5H�Q�èJ��C����e���}ک�:>��#)���Q�,�< ��#u��C��fҫ���2�kV�a�����R0hUr�Y��k�v�ʁ�ݰ�"m
*�L#=p���O��s��\�����߭����KUs�ڗ؊�q�m��(�fae&I/T/� �/�c�@���pj�y����1�$E^.��\�(���d��p�<�c�J�ZW��TP�@v�!{���)xޠЭ�v��i����Z�sv�m�p���'ruQ�m���bp�>}^�����wp������P8�0��b��}�0'���oN��̫��|�kE�nd��uj��!q4�� ��W7�Q~���Mv����[���u�K���˧�N�f
�i	�H�'�yJS����YH�?�$ tpd5=�� ����E繾I�g��K���o���R���5 �C�!v�"g2"��`� ��WfK0��=�x���jJ���)<OM"ğ�lj�o��Y�N4;�W��4�����UfNy�/�TWTc��K��`l���CR�N��ˋ̊�-Z�g��p�Y�'�;n���Fl{���	�znPZ=�f���Y�V~���Ekcf�4Q��kW��������_4y=�L�sǮy�uo�����'#j ��p�%L�
M�^�7�QJGEo� 7P�У��1�n�k^�M>�'�{�ȗQ��sbBS������t.��j�}?wQa��(قжok�Rʗ��Z����+���H�4���1�`n�\���>�sM��4��Y�r�!=x�G_*	��-�����@��TԐ����$6��;�*P�S>Z�8>���*k�Ý����˸�zO�4������Feb�A�v��q]	g�~��](^�C���d�4��6�Eo��b���D��E��db!�t������(�����L$�~�q��5�1ؔY�a^��& �a�U #4�7XǤ Qx���`i�8��(�u�)!6{ߞ}: �%�ɂ'�� �z�^�+q���<��ۄk8��;��èoaJ�*�J-���O�ڶr|&u�=�����NlQ�G��P���;a\s9}��VH��Wڏ~�V��N�۔�vj=���m�7��4P��_����h�"�����td��\���h���Yе9��>����Fw��8��%���}������`gl����%��s[���n�EN�k��/�PG���l�a���6w�9�T��<:G�}g����	���m���k�nv��h�/�-��R������F�ƥ�����G���-��fr�hL{�\�{�5	���T�'D���\Q�t!�PL�H���SQb��6�̟��BKϮ��{��{����"ow��DoH�f�*NP��H����m\�����(+.CJل ��A�e�Trp�H�O�6�05/X�:�Cʒnc?���lp5����\Gs ���c{w����z��%��f�a��ۏ���d"\�v-�NQ�i�j
������Q'Ak2��"��J�}��Q\��k@�����7n×X�@sg�z����Pgj*yQ
�+�W1����(�\��3'f3,<�����!�����|T��Y�~��$��a�G�Ϯ��fk�Je�����1���������wNO	u�x	
���Ĝ������H��S$�@���R��#�UIt�Y��5Ґ�ߣ�GB.)�=�L�&K߹��R*��1��oO=<�-x�픆�����[��ҳ�ȕ�$���	5�]s�,%���z?��MҀ��,��Z�2K%-���J�txi��;������xK_z��?0c�1��ڕ��)E)B�-.�Kp*�[g��7@�oF%�̲�����W�DEC4�,�
z3��B_��;z���)Ĕ�i�l��¥���r�I{�[��}Ok����0o�4���Ԧb��
:?n���tB0e�O�e)�g�:�U��_|��y��� ;q�8�Ɠ�����W~�ͤ�\��1����z���aP`�](��q�̀j�qH|j�����J9��9�3���JF}�����������Ĭ�b7���0c�y_.��O|Rm�`�p�}�b��K��ֵ�����$=k�|H���ѫ��o-Ã���\7���,�~z��q��g�!��d�H�/I��?��L�a�s�"���ڎ�:e�E�,��w/�>ՃX��=@��(E6�d�a*��)�� �b̾		 � ƩZ������ę�����u>��VT�Gi3��!N���D����lH�L�7����Nν�B��(p�ϝ�=ȵ,�$�՗on�V�
���4J:�Fp�ԲW��6���u:�=e��ϵ�b�0��[��t�ۇh�<�(A��ՙ,��QHx���˱cC%CQ��V��O�̉1��!}����A5�B�56w�yz	M3�bHk2�uU�۰߶`my�2��ev�K�݌@tͳ��}L}�X������A%8u(�+#�c���QԽ���=6e^ĹP�Rm惀�.[9to�H��r��_58�vςf�0(�c�������}=<��BB/%�*���d[�q�,I�	B�٠����;�Bf]�y�]���QU �OD�Y�N���8"n�֎99�<�IC��;�O��+��#|�=j�����7²��������tM*�*�䎦
�O�l�����M��J.M1�K��gނ�����\N����;67���f�M������R�7j���fk�rK}�( ��=�Q�}0=���n�Q��I5�x��� ٣��.ʕ�Gf����!tyԾez%c0��n��&	�W�e��I�?�)׬�>�U��ĳЪ���]��!d&�@s�A��S�pȇ'W�.�}j=���5x$E_Ϡ��zF��$�M�.��5d_B�~��t��$W��:��*�a
��0�Xn�M��uH��;4�ù@��ݚ�$�q��шZe� p�L�|դ_ݰ����&sU�!���j}�HE���qj�)ܻ;憹�5�&}A�R�~[_�Kv�Pܬ���p_�[�G���J�ړ�r/�ӏɡu!��h��|�!:!'�l
�G����0js"�p/$��BX@-+P����F@��蝼��tL��7�`\lk�@�ɥ�`���+�[�p��dz�'���	p" �-_N��<q�fB��=���P��t֏���������y�F�j;�ȕ�W�Y�> �� x	Ė>�}UV���[;��zle_�Le�F[;�4�s��b�\iSJ��hGه�RL�Ed�ߥn��h�ᓧIG����P���7a��3D!�j6�_R_�D�l3^L`LϬ;y��VR|�\��E�yp�?�f�[y��5r������{��%R�᜜ǽH˲��^��}%�	�/�$�IT,3$�8�`�\�&���O�>\r5P��@/_5aL�YhDkM�JvAx *��H�U������WP����saVџ�(�L��H/9:e4'��-���c��x�L�Z�GiOS6>ǜ��b[~?,��YP���=�rx�[�n�F=�c�O�d��w���5]���R�����T�<R7��YMy�7)���y���ݯ$������DRC������lJ��IE>&~�4PTJ���z�ǻ1%('�%N����b�2�og��(�∂���
��'J�~����y��a�Ί��R�(���v%4��T�,o<��giM��.�r�0�cL�_ʽ��#���hJ��kc�
"�vOv�(�;�E����u�ӥ����R���l���z��6��J���D�٤��Hk�F� ��a̔<�%.7�n��$\�-���L��ZN~��d+�I�+�-Y5&}1Ӣ��
f���0���͓��@Er6J7k�-9+K杔.O�gǲ�D1Oj�p�8#M���l���_�����2C�>��qX��p�#�0. Dn@.�Y���l,��v��SLimHI�>��?a�G! ��~��f�|^(�/ذ���'G���sS�w?t�P.ʫ>�\Stí�)��#�M`ݚ:���Ü<]u��#�X��OF^�60g`�QO���X⢩����i�+���iJ�75Tc��Z�m�H��p�6@k�?�Ay{ƌ��D�:����[�*���1rF^��q�Ӯ�O������I&���7�I����R��=��A
!+����𴸥��������$�dd���,;�	"����W�6?�[�>���Wh�xN�n-/��W#�����Lw�H0��+���Pz�.-Q�⠙}���_���Nt$�ӥ7�ښ�9[1����P�&�;lw�YgE�U��Ⱥ]e=�s/�Z 
1!@�;���lҌ]�,/�N�i����U���*C��!��l����U����d�1o]{�=��:�Ei����Y�V�*T>�i̖�����*N�UFBy����y��Rv 8��Ӗҵ�ٟ�U�Y�U4�J�_2��O	��i��X�������n����u�I�]7�N��ʷK��(�jv*�Y�9'�U�;y��k^��6�0§����4Wk�b�}���~�.<��E2�j�S�K���6�X*Q�e�	_�'t����jPDM�)X��ο��"� @�`�������O6&�L�Vt)�.�۩������>�h�;v��]���g���;��!��q7UBR��=�r�)�Ϲ�gl�q|x�iQ�82���{���w4��g� �rA�A�k]��a]�� �)5�>p����:���Kȵt����sW1�`��?,b;PmX���UP��ύ�	�����ā���y�w:�"�&@����fs��N�N��L�q���O�ͳ1�km7�abմw��Oa0,�<���77b-�aҜW��!��NQ��I\�0PW?��kd��5ۚPl~��g6��<n�G��,ϙ �SY8�
�[�wkަU� 5:Ѹm�B�S���]B��L�:0�(I*EG*1DE�4w߀�T�}b�y�1�-SeV%*ұ�_�u�Kym������}��TU{��-Oe1·\
J�7�8Đ�M/��!h����ؿ��
�ݥQ]F�u��H�؉5���V��?��*y�/w������,B��S׾��0ؔ��}۾!��C�l��*���01a�4�ʅD����?��M!C޼�e�o���,G��M�0����>�y����buS�'���=e�S����Ú��f�j'��vح��c|B[�T|3^�g~]�H�/qv�Tf;h4���vv\W"BOF"��N���uo������S��D����ETs˷�ԫ�'K��-5���I��ƅχ�|�lN�/G�t��T�������ճ2S{�j#
�LOM'#����}�����6V��-�+Z���)�퍾?�B�R (k{=*��bm֣;)=�������r4��RU$��K���@ъ��e�7�bҨw.%����3�=S�s�N�I��m� =��8�<�f>
o ���|���4�<Q�;~��>aK����aQǱx2dM�
-�2Ryэy�$�;ٕ�;O�����y��6��c��V/�?ĝ �ϭl��oΩ7��/�'j0�P�sq�8ĥ/!�v��ԃ8~Q��X�(����D��r�!��Bދd�;�]�2�Ԋ����ԓ��B.��r��@�~^����6�����8�@��KڷFIZ��XUX�m�\ ��@7�H�i��&���"�=ץ��1Y�J�0�D������3���˄��-�D�o��&�m/ �hH$5�I̎����M#��+w|5(an�X��mÌ�b|i&����i�W��y�!b&ssSk�Y�E#�pm���ت��E�\�����u���蝥�IjO�����������`jrV\��}����o�?��'�u�n��N�$�����n����t�W��+Dg�'�5���w�0���+a�>����o�{���J[�P�.�h�ےB���{nb�
"�C��n��b�������E��<d%��յ�� �VR�֗�Q�׷|�k��j����O�$�e��oҙ�Q�ǅ6<���`xQ*݌k�v�vi��
8D��U�ɚ9d�M��JH�06�~'������^�K!���� ܆���F�o�;�?�V�_ b�;(�wǣ�b���ֺ_c�Jmub��TB��
Y5�$�5GN�x.��i��(����1@������є��Q.ԝ�Yo��D�s�wB���. �Q���Ϝ���\N���k�u'��<�3�el�*���L¶�ĉD+�
�.����pm�����]e��:e�荰���_2��YT�35z'��;Xz�tn�=}���cʠmC��~+UE��}�A;�F,I�/�
��=��;�,�K�]�)'��A�e[^�1!��:*��04Q���L�F �G�>�h~s��^Ϊ��\_Z���DX�����8Ά�?k#��������:��y�{b����4�3!�6u��+�R:������F��[� ��.jTHAWޝ⸶Z/����8�`l.<��ȃJ+nMK�#Zʻ`Je������|0��kT4iv�S��Q�n��%�e�>���X��b�3Nc�_����RO�;�}��(A�&Ȇ�pӳ(�	�`��Gu$z�ڇ�~��spLN*〸u�`m�T�o>>��p�IJ��}?^H���a���±̦�\; ���/��'4ؒ"@����|�Y���&T��v�MV�+����I`�l涘�:c��KJ�T��s�����<���/�9>� ��e��.����[$���pܼ(��/y��A�tzw��M� h�c-�V�Y����>tz�]K�OT-���(p��y$2��
���@��aUF��3 /�Tݗ����d���x���yS@�
�
�b*���u�9�v꿹�#{�5�6q!�~R(S��k:��q{�Do�C)9�
.\qj�R�M����dwOkŕb�˿#*��#���bO*}�����,\}!�� 6�ݲ�Vlg��Ođ����%k�j*��<��^iN��gA"?s;�����<ư���Y>���~	J���巢dY�N�~"��񵪾���7��M6��2+"1��NlC�8��A�󟫖�4�MY�4{�����=�Ф�ޟ�4l�[Q���N@p��ۇF���)u���7�I�e��D��&��uX�,3"���K�����fDN��.�P؝֒񘓍�If/ULe!���hr,!�{�����HL��Ґޟ���B�u�l�\����yp�΢����HVO?�N���882/0ټ��3�F�4Pu�?�k�le�m��5������Q�=o�5��E:ƬDT%艺j��Z	�A+B'�4G}b{�
m�+'���57 ��	����amܴ\7��Nގc��$t
�2�ط�n�,yΚ���:�����.ۑ�t�O@��9���$}\&��>�a���(�<4r����JpR��V$�ē���i����a��d(u���"����~�=��g9���z:4�9�g����̡z鉦��6�����_��S�Cl۹��Lg��D2��* �p��2}�������L���ь�kV��*��~摆�5�k�=����d��@�lm�ԑٟ��Dm
Knn��դ� ����[`� ί��s������?�R6� c2P�gK"2	;���?X��u4-uR����,�Si�ɟh���z����(P�[��j�Hbc`�w>�v��;�S�2��ӱ:O�_��f58)tK�Gh���6��E`�AP~��Ŏ6ۗaq�	Y�8ka���)�U�M�nT�
^��N�.���
{�:��q0�4�\U�XQm���LG�F9Fl����,��~N{�Ы;4�*�]���t��VQ�ÍOq'� 8�g���NkP�[3GSB���?�����?��(�觥�������h�� -���s��k�:`��kQ���BP.�}�f5TY�}�U�G�d�IM�]���M���54�.,� �M����6�`��ޔ�Ꮎ�.&�q9JSD0t:-.	Н'da��wTҶ����{��!�S5+E���`|\���#��$I���F��4l`� �G�"�?X��m�	@�`V �d4soY���Di�õ
h���׋/��ފc��9��8��~`w�؇�*1�:���G�9PF�7��16㖫�KG$R�#�@}��1��	{X�y3;E\1�#�Ϻ{s<��t���a�&g ��i* ��TT8E�!뾎hg�1C�wI�� ��UӤz��|�eR�*`�?���d�1,Q.]�^x䭝����=Php�u���(��ird��C��ȴ�>����l>�[��C�:���P1�X��U咇�GT��|���� ��J_��NRF��,�Y^N����#�,t �`���|�LU;���IEi�� �����de/���.�z��}�X���Ͷ:�sX� �xB�:Ã�CT&_�24Q�P2ff�e`u2]����pa���πN�j�t����ȓ������G���ƣe�$�~�-X��mą�f�!�Ǒ�ax��c�i�h�n�5�u�@!�?��I_�������	 ����[i:�m�vy"��v��aS��^�Q&��{��Ԥ�W����m�>�-���5�$%��^7y5��@I�_Y����X�Ɋ*���z6�T��x�$G�=l6L�T��`ӛ��?���Օ�������~.+�u"R������S|$�h�b�kg(B7 	�����&|���D�'\{����W������-#���pd�5}Md\A��({Uj���������ݩ�����J�m�^s��*����*�
n-��JqZ�P���qE��3�GfȤP��{ğV]�A	��ǌ�Q���N�~�_b����2��&w���~�e�Y�E��Ͼ����d(,�O���.�uT��o��j�J�m;�<�sq@�7�>��d�u�y��w�Y+�h�h|�҄�;i@��ROztu�X�Y/(�F�]�iB8!���)|���ؒ��@¶Ϟ��*USУ�/D�1�{4�P��~�O�����;�Ǿ�H�8V�����+B��#���$��-�����4��j��q�$�˵�˼�t����䰙c��92x̸��j��k8�zn�_O�1A���T�`,�ڜe�ڋ��A�P���<�(����<��ΠE2�'�xt��|��:��C�2G=,�]���C*�a�z��˄I=Ĥ��S�5Kv�}��t���_��m<<��u�	�Ԑ��^�Q�K�!WF ���˷������G�$�aq�N�^s����SЊǕ�`���Z�WB��?�"=��u\��N��r!�e�8�U]��1��i
��.��冡ҾR-2��--�c�!����nv�Jq"ftqd8�R-��:�,���F�C��$����x�iA������ /�v#��m`�R���<�!=�FTPݺ����������/aÉ�ۺU�ʵ2�Y�e�׌�Ύv����:�۵�dVn� �*z��9[��h(-A���y�>���<F\�1Md��v#��3t��\� !�+J&���*��<%����U9���$M0lE!S*����rM-����W��T֏��N�������`��d��hJ�z0;�"��V_�QIX�/��D�'���Ȧ�gV{nʍ���L��]	��*>S���6�" 88?�:kS�Om걭!O�B��i*\J�5/;w*�sĥ�-�.�R�a%	Np���8yP"­≖�_+�P��.*+�����
ˎ�gJ
��+���v�ǚ� a��C��b�p�Z��8)4��Ju��,+��vA��ȁ1�0������ ���3B�m76`�cџ��е+���K��k9�?�w����2��lr��L&6hnz,�#�On��������%3M��T.������v'7����p��{�(���QAa�I���*����_D�
�ߎ3�9�>u�6�CT�0�hUI�Aп�����1�����E:'�\�#�2T@MTR�e.e�^#<Uy�}�pf)ea��1���D���ChEN�l~�lB�1r��k!E�����D�-˹3�ĥ{�`ZX�W{gEZ`[<�,K;TݝX���Rq��Bpm�Ox��f���ז�!�_[_�&�>�W{~xt��N] OFfS��N��K�jw���D�-K�����͎-�tk��v��$mQ�
a^���[�ܦN�pt흒P��Ζ.��!�$!>�����|"�����j�0��5ˉ�t��3�x��o!OZ�bx�T|�xqTݹ
�W�����iz�D3��0�{�^�y�$mU�Rol�X-�Y���,�iW��mL-${K�p�;���Ww�X�{�I�����y�P����C�<�	��iE]G��Z���M�Iz<jȘI���t ��|l�PRO��,�6��˓I4#��n��x\-8o6���H�_��q�3�u����c��oCW�A�v��b.CWI�/�j�~�Ϥ@/�3i��Quw5�#��#�ͯ'�g(�:�86�H�8�$ۆ�`P�>�q�+|�Y�iT�̰y�z�:ҁB���!��1|���jRs�M*Xp���d�X�������u�G��(<Cr�A�$���#�㠟}�1` �խ�BO�i��Р���z��e�P?�7���2�a���!���F�_Eg�#5��w�fyIM�H#'����d�� mt|_7�B�����t`Ip��M��ʶ���W �E��&\C���ɭd1P]�M"�ɘ�̕���	�K�ɓ:;h���|qT��������/�zr�m�n����G�(`4PO��W�#��g��QM���uw�.B�%B�F�f���Q�k���4g��19P�]�)9�
p�~����V6I�1��;0�m�oX���0f��N���I�ZCfa���RX���nc��X���~��X��,\�33w��Kn��#� O���=	���� �h��T}�@O�,o���_���yѡ����m��hŪC&:���ƌ��l��tm�L�h�F���JE*�Q��v%[�f�aq��J��}������By!�r�}D�[� ��Gw����4�|��o�5:�!� p��m��%W��R���WM����!tniX�v��]W���&�ˬ���9�Z���N��RC����Ǝ�6R�	����_~�kLy�=r���!�9��k��8��K,yA��ܠe76E�m3~�c>��������� `g�(��Jc,��K��)=Q�25m
]�z@�
��O�S�B�-���1z_S��:�dLQ��f&�Ѫ��{K���OE[n6�aJ��MP����<��!2e6�Uea��>i��̛
�M|��� n���1*t�ȳ<�qe����Z��3	l��0�<\�󌰓���X#2pw�5��j2m������2��l���ك����y>�d��l��/pN
�|]�����eBS�CG1s��S�K>N�hCI�tx�ఏ_a��*�۰��,M�⍜�D�s�Q��֋�k�hx�ה'��.̛�q�_I�~��exQ���z�JT��N����-螝�y25��jH���m�,"=����4� ��)~�Z̦Wr�S$�:w��XNU0 XzP�%�m|ef����݇Q��B��W��h���p�>�P�c����ּ轰�gZ|Z m3\���Y��>�C��&�5�ㅝ�K�]Cc�6��q�^XY�kZ�M��1 p�r��|�V哥T4D�+�N�=�g�U/��Ą��J�u
��8$T\��l����#9uv��v�>�v$3���i�"�`|di7}�R0*Ł��G�SAY�R6�@�+��B����>�3�0XYyU��$L�	�p�?��H�N%1+���?���D�u��V�qA�X����^q�D���I�9�I���xSk�["ۘ�����O��TY�v����#���*H�ೞ���3�U�2��ĄBA��>��2j�3���#��I疴ם))�6ԟ�O�_AfN#-�+�`:B�˸>�1��O�lM{{h���n�M-�?G� �ܨ-ydb�Ŏ����	R�Yy�k��?�$��cWL .ԕ\`�/nL|Ya�]kV�����^��Bq��:�J�d/�,��q�x	��$!�:R˃�2�d��S#���Vy�M!�7$�+R�]����٘TyJ)4�@�몉G??D�A�T*�xLEр㜐m�X�]��#Q�ŔL�f`�j��=����3a�g�K0tN����l4�h��ĺ�σo"��B�Qd�Vl�m�'�$���)!��Z����ZG����N�_����7��Җ���$ZH�-d'Y3	^G��u
��c��0a�Ώ��o����^M�]��d�c�fDmg ��t�����Q������5�R��^�b56�-4�BO�WD!���as[�I�R���p D:H�e�1$��i��������	�KWB��ۧ��6�L�?�"/&Wص�v.��ĝ	)���*�29ٷ���yeAڴ�"7GيfW���og"��y��ܟ�y�%˛�� ��Ƹ�ܬ��|��vȧ��]�Q����x<^W0���g*�M#7�Hg��Z��NsIƦ, ]�~�n>�L�X�|�u7�tb�3 [���{>h���ʴ�(���q\BX���]aQ~.��Z��=���\��־-�w4��J8t��SX�  �L����^\������N#���^�J�W���P�0mki����K{��`)�����#����d�"�8��7F�6��G����A�Ƞ�ޯ@ӽ}b���%7����[H۴p�K��.<�x�*���P����B�:Cݝ�WY���߄�ba'�bD�ͮ��g�J�Z&��0&�z�!f��<2}i5��x��'^v�!ב/J:!F�1�_3h���IL�@{�e��<���Z�YDۑ��������,���p��Ĝ�'qޖ�1���'sI���u���ļ�0b�`;@�t
�/��5s_��c"'� �z3��&�@Ex�t/���9�\P�/tk����9�q}����b��b��߶��W�W�r%�wp�5-j���7IbI���Ɠ�6����o��X�E�Ż\f�^"�(2���1�~>�` n��IH{־�	�=��I��٘;���wx)6��[�����#�R!|z�F=d�ؙ%BT��
��y�6te⭊���N�t1V��%���.�/�	%�:�� �k�D���':��A�(V�=��U���yŠ��p��ؼ8��|ڤ���W��F�~CI��à'��'�BGˤ)UB���GǍ��pQf�۷LQL�'�CG9a	#w-)顣.���mPX��BUV�	�'�w��r����|E�O�	�YY���s�����jL�7�0N�@4�s �8d['�HW�=�r�����T�mX���_���A��t�4��*Wт��[�ϝo�9ܰ3��T���9j�'A"�*��k#l�lo��2�x�(u��B�9��´��.���h&O��{��y�9\ 	̭{�F�#�<�nd�Zb�+pR3A�7~��$�NA���E�<���Q��Ӌ�@C䥔�U�E�r/�&�?��s�cW+�@�����4r�F��$��*�<������1���Z��,,CVT!4B�^�
f8���'S����yR�-c�ĩ����R�ϑ�>��z����q�C>C/��'��DeCGɆ1BN[�p"���ڡ��Z���]�� ��#��f8�D��*wG�r�6��@��u�<ku�@�y�
��v�tdg��$@�ώ��t�ӹ��Ʀ���8�Y&������SCBF���\��^R�H ��2M�+I�5]�B3��X��D_�%1xN�C�Ͱ�#� ��#[A�X�¹� �� �k��S���`�/`�Pu��)�8��C��ɍ�_������U�WN��T�}�?�k q�\+�Z��y���㻚�"s�9&bϧ���E���g�H7��[cRL���AI+��#n[(��ț0�s��ʸT/�z�4�V�?����P�t��v�U,�c����3��0�`�S�Ib���!w�#��0��6�����'���ܶ�o��27˷�T�� o�R@�\�ш@�ڌ?RA�����_�#��Қ��I
���^h���h�������,g�I�F��Ӛ�Q�(��O�w&�00�:"���
V��On�	��2`u�{�b�-z�\y�(K�D�<�@0��{k��U�&�f�`��uG���������~�������<,��;񛠓�^�@1$��A�� �BÑ��,�VgX)}=���ɷr� ��h�9�a2\m"�HX�=<���VK�M�X�5� �<&*5ܧ	�A8�Ce_E�q�0a^.[]�P�u�p�[��ћ���h���uR��|~ε(��ha#����0V����tB�%Δ�ϣ �$��S�yj,�6��Pªz���������$5���%zrlۯ�uu��ҷ����K-4��S;E���9�t���x	��J}���S�P�Q�v��~�+{#�V�̾��b�Ǿ��Sy��DP�BϮ��T�\@�J�3-}���q�,���"����,LJ�9o'l�(�����E��C��P���M���	i~&�&�0s+b_��6%��hZ��������}�����ZO[�03\�/��9Q��n6�rD���LO�66�JB%�c��5�|��Ix�抃,�A1�m_��*�
ok�_��y�z���#~�oŎ�<��^2������	UW`u��ga�ʅ�d���؆B��4�jrT�`�ϖ��l��l�Q6��rY�N.Y����m�٦�)��"��+ �m09�{ �n�������Y�þ���s��w�Oȿ�u	��Y�ݸn����:6���[��T��9�+*��k�m��2���P���Eq^X� �r'\'��/Z9�$��k���G����`JG��� ����Ө���FH�6�5'����W��ڑ?�����(8��Gà1e[��/{����0�R��R�5;b�{��3ٔF��������	������b��gi��dq��N�V�fy�U�c|76��;pl��>��zs��{(d�?<i�Y�*�L�����)��`;��5"Gu�D���^�3��� o.��FX�����9b憍��U����N[�E.P��F��	'�h��ڥ�"�9��SO�b��j�/3��|	$!5\�٪�H��Z���^o���9�&;볝��Ď�m�Hm��dyOj���0g��7��n"EbÐ��>S���u4'�V���%d�/:ʴ��r��A��,��U�ItI�ne�Ġ�����G>�J�°�=ci\_�1c�u�j��ˮ"y�Yٲ�J�Ŷ�[�y�����f;�B��ê���m��j���M����[�`�b9�}�����H���,b/nv�CU��>rt�ɪ来��ʹ	2D��JN��fƺ��C����΀N��]�C��r�7}W��S��9{����	��YѲ}$Q�����ב�� �	k�{_l熜~Tu79�� C���=�/�g���$����h�B�u���:�-x�M5��ԁ�^O��:M��j(�Ք��`,hG|?�8��৿�=��,c3	��jl�y�ʿ;f�,�>?t7G���IXznaC��T��ƹx�	0[�MN����\Hv�t���X��UT����a~'�ģ����:vb]��]�V@���9��/��gᶋ>E�t5��	!��J�iӋ���y�~��ĉ ��mF�\	!/8��Hb'��m��O���ڏ6.F�|��7����'��9��q�ֈ�$6��;GOòp��w0u�>�l�4���;���H�
�����x��!�ZL[�?E0��'%�.r�g2z.��~���k~Q �;��(FC�m�!�a	����³���a4�5����3�p�-��C��5N�!SϏ�c�Q~8�
L8&/Q�_��HtS ��G �Lx�s�v�ޥdq���>	���"���*�-��$	�g�]��+�M��V�:���k$+^*��[��)�|���������\m�d��Cp
_��p:�M�W��SIt<���/��b(���̘���t7U�ջڅ��;FD��sg�<)m�����,B�����EX?N �(�h���"ƒH=-��xz�w�C��-�ϕ�:N����Y6����;�ur���*����H^y��\*�_��U�΍3�k%;ԖZ��:�� �#��H�o���uG����<�_�֣=��b疲�6�	g~�)�_�e�hY.�Τ�hP�i�>؜zRgc�g�+��Q�U��"�e0ݢ��e�i5������dҾ?�8]$���A�I� ���E�P�ގ��<*U��;�$�8�H����#��D�f}AA[3�,mF׺$�l�j�fzw���u/�)�����h�ZHqA�S��"�t���ԙS�ç1,���p�@b�?'�R���n�~!3�}�C��e�^�_R���U���5i�Rx7�^��ohI�_�1T结(q𱸼2#[<���P�����՟�2!2�z��r=��vD��^��ɖ���+Sm�����%�����}��5�-�2�~y��s�����)�⭊ B�R�Mb�m�#��k��zд���G���V�̯"
7a�3��rN�"���`.�@;<(�XU?�f��V]��*��^����h��́��gp��Q����Vcc+C֡���P}�M;�aW�śBx��� ��|+=m2��a♱D�rj�\�o�w4�f��70"��H�KV���4WXG�'@����G$O2%Be��eu�����j�u)M>d�"��l����X���&#��J��_�^u�{�5�����#o��w�Q���!�B�vz>Į�����>c(+	��eB�	6:d��1K/ɭ�sy�Xo*M�
>�N�_�AN�?[���9�q��.�lB>S���s[S��* ?͔�J��O+}�s�����v\��֯���e��c氅?.�r��B��F�h�$!���9�:��	B����3�}:��qn*Ίn>����s}��,��B��jK�G�0e�}%�� Q��y��qjW+��眀��S����d%C�1���-כ�ء��D�Lc���]a(j��I:��3�G�^�m
kG��`��~����2���������">B25��I�QsdV�RC]4VJ1H^H��8I���q@a]Q'δ;i��gz{��L�х&� ƺ6��g�K0\��+塏�f��3ꀎ�{|� EG�����,g=�k���}؅j>�7,�ǎ�8������<��S]a��
��0kR�~aI�U��6^CH� ��:` /��0��rS�갇q6�]4Ss�+��v�5� � I��L?S4�o�{e8"}�<�E�I-���.��Vv1�x4\��ߣ�B�*�H�M�t�:&L��^É�m�yz�'���p� 0�}-�v{7�/�
"�+]��aG?��2�+*)]��[*�hݞ��2e�3x:��W��Gr~��uS��<����}Vt�;\
2��¡r���o���wŊMf�8�gD3�Z!^��\ Ɗ���\kH�d�U���U9��EJ�5G�D�N��e�EnAm�;䅻z���Y���#���B2iR4l:��&_S~��3)+iǝ͈�,���9���{Z�bC�8��ˡ��r���i�8�s��1.�v��j �h!��	����θ	���p>b �F�8�“�Vmψ�/lCi�1�)Q�l.�,�s\8�I[u;�9�[@1���ν�]LF�R�A"�t�%ذ��ڇn)iP�V��+�f1�bh~(�~:�$�릭�]�YE�o.j������Է�;S3�	s�֝��yHQ�����-Y��G;�R�W=�>�e��!�[RM��>����T�Cv�98x�kcw9��� ���öz���f��/*�5B�5�K�em�w*M��\8��.	�I��A`���4�=�-rz+Q!
��ü��M[ؚh���Ke�Q1��������`�ڜ[W�D�	C�)h?ؑ����
U�Sa�� �Q����s���f�U>��/]8 �K����K��Fr��Gi�B]�_nR�c�L�<�|s��J�-��RT���LhgA�lsTd[���ٶ	y����B�_�z��ug���K�} ��?,q!+�+��������I�=���T�6H�4�>�$�>�i�����9�0�Iu:MLt��7�]�w�)�Q�<�a�}�Dd$�g�N����x(��V�����0ݹ��D_�5J�̟���,���Aĳ��C�|��٬�]��g�,�>̺��:ޥD]�h��_��_�5!:�oS�˲��>�\�@SC�r�~��Su�<�Z@@�o3gXOE&��ы�p��Apt�xu����l`�p�4jq�R���Ew�|l^�5g����5v!�e�rE�[�K���UC�:�,���M;�S�1��n���vw��qƊ���v]'[��¹���[#�x���I*s?3Z�����y�~d�@�[�N�ς���2WJH������7�|d��|�`�8&.=ʟ��}�8����SO�>az�����V�u��/?��&� �P���<)"%Pg�Bů�<�V�D�D}�l{^`�\�:&ݤ�D�M�b;��E�
�{C��D�'�c���ZhQ/��u��5AV�&얘�)�-w��8\)�0��>iVQR��B��};��w���A
�?�!̣'��gV2ƚ�И���iz�Ae�|�>��E�}qTBEq �6���,��z}m= ��o��S����욝H5Zh�R��2��#}�4�U�r��e�wl�l8�c��hH��4G���ż# o9�ƣFn��<-� n�,���$$ʦ�.�	b�_߭%��yɥ́t ya�10sx�uN���!ʤ;.<Ơ�����py,�'��O�z9��pn']��>�uʙY[s{@�{�~=��s��Eml�X6��1����g�ka���]k���`4	�J2NW��&����|7�S\�������,Q5���h��(S絛Z�-�	-S,���Q�h��0��JcajsHe&X�Mg��r�l���h��P2e1��*WA�ɢ"��� ��<��c�u�n(:��k6j���_�R�	K���Ꜣ��uL��\�Ȯ��zc@���)�k1�3�XR}���(W��h!�(�.����'Y���/]�B��f��DrtF	-�+�ɯI ��I����[�y%��
�WH����xب6�TH~�-�n+݈l�p����7�Z7C�ԇ���ry,�*��.�9+��J��<(O�I�O^��gv��
~r���qf@�UB�wm"��0'QA2��4wW�;�#37�ҵ^���@�2���C�O�@`'=Kr'%����
�ad���%lA/���Z�?p|�K{6�I�BǓ,���M�$��gl�R�.�\���|��?�tH�	ЏxV��V�Z��Bo�D��N>�|�(�����H���X�N���^��T�C";��Þ��������#ܑ�VC��oH}#h~��xq�5��Q7D �hns�~p¶��~�w	G�1ҽ��{��۩$�.=��a�	3	<&�yhi#����a��(��:,��YE�*�-"؍rd����ڍA��r a��g	*��q��6|m��.�Y恦c�~�iN7�ܤ 	�_&�$���L�1Rnv�����;m_G�r;_	� �`	�e�6m)�R!���HA��l�H�Y�uS���_x%&��r�fu�����L���g����n�����3�1�=��lg 1�9N�y!**�0�8�Z)�����[�✳=��ȣ�`�ŻtV�zh���ĸL���b�T7�o���� �H�$�po �o�7�S�.�T������po�[�v��>4�M��l��ӛ�}��>�j�>_84�Laqg�#X�@%Zp�����,�~��3�pꩍB{�l���?<��^&����}�^%�@zR)$l۵O���gǗz�� J�+��{�����į_>�A��W�\.u�鵐E)?v-��Z,~e�hhx�����]>N��� R��--4i�����G/Y+
�3���x�������E�C��ZSO�(G��KE~������ֹo�ٍ��C��4�K{$+����ڌ��!�J���(@��^�-L"��)�Ge��%_A�£S�G
YQr�?�?2���h
�7h�d��G�����W���_�+hFy�������!��	J�vt��4Cv�5�PhB���$0���-��n�Z�$L[�hZ!�G{�V'�uĠ�区�-�Tq���/fT�1@fr�xdl2䐥yo��{`��l�ʟ�Xx��|���Y�|�2����&�8O���/d��ZY�- �ϯ�e9��e0����'�,�+T�ɗ�C�� P����SS��}f�£T�4��h`J�u;�r�_��skJ�(�#
*{,������ض����۪Y�uH����(+������c��Ԃ��Ry�k���k:���Q�3otN�彜�<�D؃�'�-�3@Va����^Uw�V�6����A�X�^	�L������]#�!�����V��O�|�[���hʤ/�uO� wbl��Y�cU+�D�׋'��O��# ���̖����AU���.��a�N�Ԥ~1D�	L�b�=2�����'0O� �J��_L|7��|4o?�&�Bu7�t3r�4�W���W{�!����qy���|�	��jVN���.#�P�R~JL���pv�K���Q��v^Dc0��
�L�pI��o�5�vH �Y=Q����^۔-y�l��W�S>�0bb9�0�gn����,S�Ø�^�'�L~{�@�����?�~*툱�#�0�s�Y����Rw���ҍ��ɜ�y���R�}�.����X��� �����i5�C�X�}7*d����-l��[ޮ����6(f�ҵ��wd쌶�����]y�"��[���<!��0~�X�j����Lh��i�Y�˴*�>�<f�)�n�\'��2nX�ѯ��T"[��BjО?II�g�\��y4p! ɪ�RH�tv�t߰������צ��:���j���K�m�0��ssڎѽA��A\��9�M�D��]� ]g�_�G��0�,l�����QX,����	xeH�Zd�g�&�$Ԍ��0_<=��l�˷zH��`ni$�1�����Y�P�6?���[$E����¹]������UG���m�ߵxX{X�ㇴ�)ɷx��fK�y�֠L�h�	���Z��9���Jm�~w�U��@��y-lG��a��'��m	)��\tBЬ�����g��t���lQF�_�RKb�ڋ=cV���M��;�3"�=�7�Zm�Ǹ:�|�E��#��"^�gYQ8)����R�cK�hOn�6�~y������f6kLuw�g��0`��u���З��d:ޅ0�*�ӖJf��^��P']9����r#��߷$��G�d�k�y ���@�̣	[؆q�l��TZ*�j�*_^�6��DK
)��[X��]����J�(��w����D�#Q�f�P�ۮ����z��)��������i�#|:�m�3�ښ�;�?M� ]������>0��UmL��ۍt��I�8B�68��A?��_�N�����P�W_�f�U��J�PRx�uՕ�6y��嫯�U}�`O�2��n��D#��Sv8�ttO�����"Zv\�_v��'�$@���� n�eyu�F��ü��8n_M�j�a_Լ ��̨C�����ۓ�� !6��.w͉�Og���Y���oh~o�:J�X��O�^�VF'B��o�P"V.�SHw���k���Q�N��=/*m��M��u���@|<όB^�D���������f��=�#3 |U(E��_��31Ϣ����ʥ����yz�l6�F��F����k�&��G�r��А��s�����!����b�"Tϗ������UM��[������$׿F!E@�����>l9��W�]J�|�h�?��Y��H}�l^A��d�|�W�1̀�o�K��+mІ
��Q���B+[}�*z1��-'�s�vKS;�,�4|PXQ���?_����6cMt7袡%j���}�)�#XL��|�e�I*���r�(3;�\��{��8�D1[���ؕZD�����x�1Q[~*�$K�T������oʧu�l.X� �9󤬏�}q�{�����;�D^�ȕH-����P��*H��H��?�����q^�&=	s�5�g�$�]<�\��j=�*��Ҥ��{�}6L�L���4�z�f�M�����Yg�O��AP�R{!jy>�;���ۺ�0f���d�'߉���6I�rrw�4�`Q����NI��g{��y1!K�@�����t�+s e�KA>��5�� -�@��ȭŀ����Q�j�L�BL�Yy~��iJ$u����6�qh��v�\kq��KC�i�������xC��JTՙ�Ք�Yv�QBp-cj�vY'�c꫶rd��`I��Ƿ�big&����ƆM���^��Ъwb4	V�%�����)��S�[�ǀ���G�j���Iu�=��RG��5E���>Q$� �s`1�D���"�L8[�ݓ�^������-��њ&{�ie��>�n��@;Aau.h2�_���H��T0]����������c��|�;���#4�v�����T*���P/^t]�\�cȑ���� ��GD|�R������yk����?	��g�l`�'`��Mk�\E!<	��JSA�	�*�����[w���s������1��
)�	�@:�� f���h�O�=���&uF��5���k�ٷ��:�a
�Z�=Y��7�]��	�RgΡH��,��bOi�����C�nۍ{\��q�d�<��=�4�� �M��:��~� FF�v��=�i��j�2Jjzp�u���K����]@�(�녷��lW�}���w��Ճ+�ln�7;�� �7C�7Y	F��t�)�{�+�Eަ��Ξ��,��]��=�!2��=:���=K4:$�Gs2"���V����P�\�@İ�y�Y4���M?L5��z�SX�t¢kҺ�z�F��x�#�$dU�<�>��vL?�38KMt
&�K�����ݤ�Ҡx��H�=��-	�u~�뿤�ӣW[���7~���Ռ�ţ��3�\�k&�@������K]X��o��&�Q��v�vmي��҆O����ӳd�2Dj�Ϝ��IE�x\�@�9�Dx~���|��Ht9�P�2�읦�cU&p���/�De}��B���x����4���R���g��Ϊ0�+;���8&ւ���G�828�/w�X�.6E�vy�*7�ZL���u&-�	��ik��!�}�)N��Ow`�f3:�l��L���3:Ĺٻ�֨�ޘA�P��������H�1�Z���mJ~��_g��t+F�"q�T��i7�N|�[P�O�H )��{��'?��d5Ti����I���]�`�/-��|������������ӵ�=�"s]?���>gqO[��.sƬ���:�����$��ɾNd���f�+_h�n:Ў�� T�R����'����N)|ܢ�t'�1���6��-�t (\9�,��pB¾�ϙL��&�X���>���9K�����] /�˚�㫵�b��ɱ���q��c�{MJ���F�amN3Э(��޾�/t��XыE���|�ծ���%.q����1س����z��	)eٵj��w)!�* �Xv��{��)�&T(1���NG�Wh�!6���y���	~B �؁#$�淃l9g�<�r*V-%�Y�<Y�6Ì�~�f�w�3�ꈱX�J�J
� ����{��~3�RF�����7A�5�	��wJ���?�*vJ����^��%���&�$_rƣ�Ӏ����K���Ҵ\3�22ſ��α��Y\����`l`�� ���1��_"XW�粠^�~��mLJ�j�������@=���jk���lsT���}��b�G�6�~�)	ո`.�,��/=�i�Z�6 װWV�E@���նO��s�o��H�P��j��Ķ"���a[h���&Y����7���3RI��Õ7 kǨ�\�$�Og�A��"��?:�gz�ޑR��Z�ש�	��弳!$YO��c��W����KH�+�Lc J��'o�B�G�RLb�͸����	Ҡ��Ǿ�U�ĀH8��s&���pj�߾����٪�C`���|�d�Kh[�Ľ�XcPb��GIh���_��0�ฏ�Չ�FoCF��*
�aJG�Gm�"0��MH@:d���sNg���r��ᴂP�J8g>ȱ��;!������z��{c�;6篍+}����F��k��a��cjGߝ���IA-3cM[�惸-q��2f�^.���i�r�d��R�s�������N���)�S�&�8P�k*�Q�t�xz#^��vh���޲a�D�v��������=O�@��Em{�I#	�5�"s��A-���Vi�	�Z��䬃���l?	�Uޤ3������n����eʦE��-�����<��z�3o��8�x��<U�<h_ȡ����OJ����R�{w
k�̂--�"���[/�k�xAKc���e��@��7w�[}d�热|B�_i-���I���v'д.>;Cf���owuN-߲S0Xzq�����G�7̀p��YWV�v�ab1�����Ζ��@��6��IgQ~C�#8�����ڝ�Z��?��{�n���?�<��[h���롯��'|޲��z��2��15ֻ5��<� �
e�ac�P1\Y���;1���H�p��� �Z$	�Z�w�X�tt��� 6#���m��� ��e����3EKup����O�_ �W �B�@�6��\܉F���WC�g��V�Ic�S�n��r?)�0����>ܸ��4��@n�T�t��|����͘�;ئ���p
�G��OV{H�G��@_� �>Ө/$Ȕ���ζ/n^k��6x�]��g$'a�R�YP L�Ь��QS7���ﾗ�1�Fe`�lf6N�4�4ΦΣ�wG1��,�m�$��Ix6�d)��,�j�u�B�^����K� $|��q%[{7xYF�Eݕe�-�r�t�� ~V��;N�Đ^�w������?��\u@)��;���:�L�kC篋
��C�AÎ� \�G&�%tk��VO��n=c��.��=�8w�t���Y�;?��	d,�Ŭg��l�.�sP~�y#�c�>�jC���J��s޴���� n\f	�t��cYՐ���^�0�d����'�aa2Ŵ4Y:��	˦�f��-b9��S���rԬ��B�Ub�8�^ٟ,��u_�Ȯ�N>�G�l-[��6�!S����`]O'e=��Wc�#@P�M	���τ��ȍ���=:+�B����fE�˨����p+�Z���]�x�]9�8L	 vVp]/��D�WW~�=��28 ���#	%�NqNZDN�lǠp^� d��I[������|��cL���tn�7���x\�7�?���U����3��/.��a��[F���h���W�2��]���(���1���ą�c9��	���[9�y$�np���f���f:�m����k�@`�];W��Rq0�XT]��䉮�O��+�4�~|������ل.l/���C�g�����5��9��Oh5���@�p����.Bx�U9]���L{U�M҃\S��j�,���-��"�Ǽ�w_�䆇�*�EHF��2�L�Y@�{n����
��M��P�Y�⺅�	�%? ��u�6�1�k�Bx�*]д����]�9O_��u����`��i�U�%}�㦢��Ĺç�u��ƾ��>��ƃ�YC�� =Y����"㔪�:��$5���u�+����',RAw�_�)+�XHh�Tg|xO������� 
4�����b37VO�8��Ar��ꎏɊL��l�-�
B-�$踋z( ?[�G����Nf;#1�z�i>���F�%��)_$pn�x]fR�A��n��&�<bP�Q�~�:��W���%c*?�2;�$�n«U�P�_���b�  qd2�zj����V�5Z��)���cg�k=�;�����2uH5��M�f�8H��]��xf�}���DV��?�p�bh m!���6'sB�r����#2�j�ė��j��R�]e��}��Ÿ�/����ӂ	=�ƿ�!�Re�z꩏���=	I�Nu�nY�%����2���C�Q�D�����k� ���P����C�N}v^�HЙ2�hWo�LZcW�&8/�E��5�f�pW*�rAo�֜E�Er�����]⚂X֝M�F�ʞJ�O�H��sU�� OL9��w�_�
��MضL�O��VV��9sh��~p>��Hd1�����)����^e���_$Y�^��vEijέc<�u���(t때w��<��+[���0.h�9�{�F�'�'ƳG&
��,�=���̅��k�t��K�m�Aq�����hr��KCS���R�uУ��!��W�ɒOr��,�����a��K_Ȯ�~X��(|����ƅ#9kL^C�.���uo��p\r]�9T�+��2W���lG�Gڥ�ov��e<�l3LZ����ӗ��)����ѧ��\ٟ�ث�~Sݩ���d��b�sU�,.�h��G�!�ު E����+.d�'2��:���/Ztj�!M�G��Ҵ��b��~�-����s5'n��+R�b�ͻ�=U��vg���هs@����&�˽��i�޽�&����(���9����uԠ�+�qЉ�[5;^Q����;�߾>MԐ1�uV?Ī=lD��w��Om��Hl�z(wp���BG���!�{ٻ�VZ�o����q�e�ܒ�S�3��IJ���0زc�X�x�ƃgY$�@&��X;�ZT����d1����)���d�Ư�A��d-�c�Jgr̜:u =�}��Ѡ����O��x7�L���\�mzRj�z�A��l���G��b���Ͳ�oT7p/��ݏ�|�O�F(�)}f]s$�۳F,n�.�4�s��d=8�l����n���)�̃@4����"��^m�M��p\B6�V�;�~Fgs��vB�I~�V̄-�ʡ�TbQiZ]9s �IOև��%U��(��7ܶ&�I=@Tmf�����3b�����s��)Xn��*ڶU<#�C�Ol��absj5�O>} ڬz���Io����OL�$�҃]�×��]���M��Wuߐ�1��&%	q:�L�f�U�?��J"+�����;pP�6\):�J�Ww���n2��:1y��%:���-�5�\��A���PM�'���Mj�7�I�E���ۜ��8�8����C:ڰ<a�:�G4���N�V�|8_qҡ��ӳ9՟GTL�8���v�����?���������6ח��H ��ߋ�Yc4|#3qbة`��F}���%��^�*��_��n���	�����	G�+�!���C�)!�0{�Q����Iʑ�m-��yr�?�o2��~����H�;˒�f�v���%_K��Ѹ#p�#��=%���p�R�Ca��h'El~�=K���|�p3�+�0;����,g`#�X4Z"WS��>ql;�^/��1@s�\����pc��H%"��2�Ǆ�[k&)І�*���ƛ_!�3��o@����A��&~��괵�������Y���a~�}i ����OG�NM��'�q��:�!Ua(y����b� B2u7�6��':�u3����e{8�95��@f�g��Ԙ�D	���V�HC�̺�I��^����D�il�9˶�%{�F�)���JM�:�OD��a�u���֦���0#��.��X�&&tI�k�b!aTA�*���#o᫆�V� �ZI�@�E��w�2��U�lg�	 �a�����8O�x=>��ə��4��/�|��c}�����t�G�����Vϑ�'� ����'V4y���ܽ�륮�� �Sy�%�e�h�k�na�[/���C�s�͖Xf��~O����K�Ɂ�`ӣJe�<e��L �9��"��@:������X5����2�E��ء(=�$����u~I����^H`�2���`��$�
_��Qt�X;cX �r��ٝi���#�vmY�B�?Go�|��fZ��NͩC�@�4�&�A�'g���A`?`K>	^D&�WM�A�\gy3Xd$�9
ٟ�b�$��Ϯ���ɞ�V�M ��6��#vF�k�n�$gae"������˨7��f�U�G�\*�B!l�o��q//�8������� ���o�6�K��7S��N̛��+�9� ��#s`ɞ�;��-;W����~�ρf������#� Z��
�?t�̾v�g-aT	�t�+J�H�ā(�ð�=�l�eSH{��N[��J����R�?%{T��X[���'N�<���s���P�ޥ\��i`j���?�U1Bh�%����u6a��N ��v�H:ͅghb��uܱrN��T��E`=l÷��=`dֵ��?84��Uě�����<�k�1�o��&~`����et�@^�kb���pW� ,�z�� Zp��pz�ꐦZ
��R�!�J�Z!���	��ٻ��_����4��X,����2U9M�g_H�:����)r$����İ�5̱�BN�(�ܷ�̅�u>��m��5�`��
�(�6Z��%���,�d�n�vU����~,�m?f=��xn����0F���ʶ�/3tگ��Dl�у���.�{:U_�����|"g U���J��;�kOou�G��<�M"�(R�`U s�����4��w�kf�%�Պ�2�����#�z~��nG�؟����	y�s�y0�o^54m��3yw)�����&�0���h�V����zܠl����bNP^��1�ٴ�x�����vc7O=r�o��W��ΩqN$��ٲ� y�X#b��?��ΰ��!1�R���~ؖ��}�S��b���h��/K���8����U�Ƚ²�AɽrY��w�l3c+�V��_Q����_��6O�����&S�ܸ)�������o'�����q��~H�zɚVy7'A��9h$p�h��a ��/Y���b�TV��-[��ݜ��������1j0��{�����a��[�c5���
�Μjr����k_R�i*W������{F���8&[va�r��x����"�PY��Y ߒ&��es�z�7��]^q}#����
8�֕SgM�T� ذ�dG|�vC`��C[��U��:4�h��G{�i��'�O�}�r�2�}��ֿ6�,c� ��L�G���קB�������CB[@P�1�&d�OHk�Oy %�dِ�Q��Ec�~�[n?�-"��J���g���"z8o���궑�P/�\��InFf���k�x�P�l��G�M���AS���&�O:�`V
��zL�6�k@�.ATz�z�q�"��䕻����ÝX�~p: �?��]M��%{#��̓~+>��㺸m�7r'p#��,�^
�÷\��|Z�:�y%(��ɛ�)�\'��I�cN�yYg��y>�N����sW+�%�7�A���y�`T��Az bMN�2���h`�v�&��ѳz�r����9���Ɖ��x�}�"?Q��]$���e�Q8�%���"�����T��Q�bP}>�u5�:�f�lQ\�����Z-���x��a�����d_���n&����4�Q���H�����Ҍ·�y��ҩ1����`�+����/�&P�}�-�G�2�Q��Ѩm,2-<�Qxm�^8�d51K����YEE�����,)����sU�m�i������w6���C����<�3ǘ����mJ,�$�b3��߻�K��2"�9���c	� �?���S��2
��[��U�;��?R��m?��9�Δ���+ٕ�;�>�P �mӠ@+V����C5G��_��e� �?�D�����Н\sM+�=��f �YQ�5E�Ԩ��T�	��S�Z&󃤝�k�U�yM!�g�����+��,֦ z\��vOi��Exv��_7����f9��L��q�ȃ�=�r�HW����E8�~����V��~1���5��m���I�OJ�bx���䉜-��i`7T�v-�e�������7�t,ñ�^F*��Ws��*a���#)O7N�[�u!� ןdٸ�}ɾ_��L�*��C�}����'�.g)5�5І<�m��@%D^�؊$\/��r�o�	0A��bZ��9ڴ��M-/J�F����PG��#����׳�kl��� e,+�v^Py�_.>��3�y�ZA��3�܍�s9��&���&-hvě���v���y��9�21r˞Ӿj�Q}�ZR�+���C�������AMj�	��X��Gn�m��gc]�ׯdԖ|ڣ�&NN�j؅�"�ۧ`$,M����.�\��� ]N�^��>/+`9�q�u诞���n�;��Z���n[�_`�e�/g�x(=�EW�J��<��	�h4���7��3)�=�;���7�m}T�'��u����C,/����w'Q)�<|��@"�@��h�t��"�Kq:�

����>3����i.y�l�7kC/��ù��<Px�S���̳wf��Q,4p�_po�z��{�'B�$		<�V��c"DI����Z����!�xt�Qb�y���$�G�0�_v�jGqZ�K�@�#��J&�Ϡ��O _u�ni�æ�x�#)�/�K:�8�}қT�ԙ���4��y��·��s���c~��/u|q=�D$�nb� #��X�1¶����v���v{��X��������].�c�N�N�0�EҨ�\I�A�O	 ���;��Yn%�� "�"Q����]�g��8��
�y��UE�������'��v���5�ǲ��»���o�mI��G�2�w��c�}3le�QI�3��YrT-ZjO�rf?�u�a%���X^nC�����wbm� �Ԟ3&)X���G�H�����������$��ձ��n�dR�2?����fmyj���lI*3�h��Y���� U'N꤁:n�]�6���j�Ex�O���G������v�
�_Hd4�J8K��Z�'��|��S��iEʞ��]O'�qg���m�[�G�lӞ�~�9' 4.l�@�
.�?�w�:��5(=�������L\���Ҷ�3��BYy����\�a���݉�*Jr"Wa���F7[q�`����n =c�c���in!�n��eɾw��:�H��n���!&�""��J>3��em�c���k��^MO��۟�|�>�	�|��e�w�;?&߇�6VR���Ɵ<q�J�~�Ȁ��P\+��/Oz��=L�8�H�\��L�M"�5�20�
�}�Q9���P�
�W!/9���D~Rp��@���%[֭���S���Ҡ7���B�	�eт���ݏc�w#��Q�*ܳ��J,����w��gDM,������Lm1����9C&�w������{�����f��1�}�LX]�;��ҋJ���ّ!�e�_C�a&`.���q����ko)?`(�)�щc��2��	��Z0<X�R�7�����.G�r�7�tE��6!��S!5��k��-bw�e�y�S�|������d��}%��g����m��*��g����|�~��dK<�K��H��
G����4ի�&�tH�NbM�j)���&*���ؠ�	V�VF%�s����4�y�*OKN�w�T@m�	��w�`��v0A,����iZ���mHɺ�E����a�8��˯_^��f���T�\8C,ul�*lM���1�"�
#����Q.�@/�,Pm����Sy��YFw�Ё�>�x�-*>&{�gz_�����/\��]a��U�E��h��,`�����"�^�<]�8��A��;�_�§���g�J��`����E�,��)�H���7o9�<�*�|h��|�Z��q�|�����[a酞/�o"e����ymhD��u����Y���dJ���kp�(m���k%d��9Z����˖r��;��C��W�	7�T�~�dF?�-��z	
�kre�"iZ�&���� �JY�w{ʁ���E	B��!p���f�Q"(�܊k�9��y2O��l�P���!�%����oe}@!H�4���A�(��� 5#��R��a�C����<A��k-ŵՅ��֬�2�C}�K��_�av�B����Z@��P�m�����������3k�S:���-���ǈ.�����3�!#v�N��t�K�����O>���!���0ð�Ћ4�S�)!�[���H� ����+�����/�v@�6e�m��K��ֹD}jt���l�G�;6�+�,�%��9��풄��`��=^p"����NC�ޖq���Ԅf`XV��Wcb�v]��b@Y�)�g��n(��l�,+�o[�(9izG!��͚���y����b�K�W ֺ�R+.�q��a���88��a�"����_��n��9UI:��I�mPY�W���҉ռ�ȼ6V�D�iM����L�U	�#)��GG;� W	��D�:K�K6k���l7��:b��!��(5��/F�s���j�|�Y�KIl�?��w�^k�}5��,Q�^�-Z�d"�A���i���
b�_�'���]�|�·MlZ�~yTϤ��3}n�)���.ݝ�l�(e�10�h��.�إe���?%�&M��n#�w_[�DZ�pv���;���y��먮��(�MpG?G�cW�I���y�������'�sXL~.l�w�X�7`��>"B-_!G�/9��K&����QsЖs���B��P�)}ܶ���Tw-Cq	Pc��A��R,�P�v�jD�]�����Xl;��B��8`%�����n�S��r.O5,i4�48�� w�;����_��!��3�y@GΆ6�
�)�\5��1���G�S�xHQol2�1,���V����g���2�+/.�8�ʓ���_�����sp�i}f��9��(�67�i��j��$��7��_��0TO�{�h���+�=��'��'Ő�]�x*(�L��*Қ���\�����Q�"�\�]jxDë���?h>�FS�u#</�����/x����=�������J���4�v'u~3�����,�A�gb6�WE���n��W����o�s*�R�X&oj搥%� �K���VBX@���Ҟ�>���2�daȬ�Xc8E�h�bO)��H:S�Ί6@�r�!q����m!`�b;���C�w�=�I]�$���:��2g׽O}S��� ����g\C�t�)Vx�j�����'q����5�!�s�p��Z_��L�y����1�B�i*���Q���CD7*��ͼ��p���AAx�0�!. J�@����G�<s�-���h�)9�Ԭ�8%��@-x�@��������F[-�~`g�mD�Ćc�rwPC�>J'���hn�Z??+��?��,	2�����E����j�DS:�$��3� �w:$5p}T����c�x�'��0�# �Q���Vs?֯���2�~_����W~�v\hR���D��}� ��?u�{��w��غ���^�~^�Lד����3��+G���v~ U�餺��C���a�"<4B�t����$�`��j���ܼ˩�u��m=�,��f��P���+�/V!ɢ��%�/�
 +�ى�6%Z��_{&p�!�K�ҥɀ�¤OH��܆���[��/�-ǝ��k~I�������H�	/A�`㚝'}�.j��ېD���������7ȼY|/�fj52��l��2��rK��ߡ8E�����Ya�*��I�!�����g��S����,8���f��P���T�c�αBgc��7��|��E2'�s�pFW�
B��d�=�Y�ь��<Z�p8�H�����5YF揭w�@H����L�{v�g�i3��{WCQ�^���F��l_��w��e�)��.�+��\Wfkui�-���,�z���6�3 ;� ���&V/L�m����b��}��G��;�/��x����U$�4)R���Ԏ�	�e���jw��tD7P?�&��\�Z�-�ʏmbl�z��k 00��B%�m�`	�e?�[n�	L��O����qa�.R��Ц6��7�su}�2���J2��ѓ�vg�!YW�����S�T�y�X/}x�[ҏM�68�}��Y�dKez���Y�����P4�l���`u�w7I)p];�<M��= n�vB�j��AeH1/�S�Vn�V�µ�l�}i���a!��%h�dۼ_���[�l0���x9�G:��>mbt��Ʈ91Q� sIC�@��Cn��Jb K��g�7D���*6�\%8�B����Ί�#R]9ж�P�F������k�&%�;����	�~�R�R�תƢ�թ� ��f��<>jNø��#�B��k�¢�h���.��l8"��.:�z�<�f2e���m�e8���<���HbѪ��1��FqU,��l����@�GL���5cm]u�ߐ�w6߳Cz�ciV§�0*1��������W��̟��jnb���tN>�^[�m����BE�E�	�lf�N�O���{��$��D*�EUsK����iXZ�0��L�1��0z����:�XƤ����iZ�����%NyP��/㾠��-̞	�щ��"릋�_?!����ןj���8�a�ǻ'A�!)�1�9�a\���$�]�4�Ld�.sRyip쁭F�M���@0��
� 6�~��|d52��M�o}�:ߊ%�*DNvx/��B5�8g��O�*�G�\w��/xL��<=�p����$YeϞ�d�@�ju}�Aa�rЈք�Iz�e\@_m�ߢ�C�&o���Iom�~�U�
ʯz��F֔5�:�p6y�"��,�ELc����Շ�N���FE�����B�aA3��K�\�
����C���-@`k90�A�e������j�8#WjY��O�Ʈ���o#A�\��˲<XJ���ɞ8O�����7�"\����	Q-�Mc �E�*��H�\��֨�n�]4q�S�eR��v����|:G&�Gi�a�at���9�1�^�v'�@I��n�� ��͙�'���~q�e�U�&�P�^c<�MN����/.C��*�d�, ɱRK(����d�Z��H��m*l�F��i]�� �o�찆H+&5�^ \���uH��]|SA���(�A�����c�IR�=�n(�%�c�6�ov8���}�+0��g@>�߲FϏ��z7US��\ye*��xJu
���?���L�O��M����T?�����h��~���j07  ���&�[2N� N%����ׇ�`��A�f�M&���bNΙ���;6��V��}��^ό�?w2����-�^𮤟��2Ld�-�,"&;Ȣ�{�V��N�26�qR̓����=<h���4a����t�|m0���v�C �-��, ~[#Ek�u&K#В��v:{�A�}�>�|���$���������z*���d���đd��&��o(�<2#��0�V������U��|%�[�dr���W`}^!+����w��%�`�!^���;���9��d9�8���-��]`HL��\-?ʰv&p�n���%�tQg�=��v)vড���]Lxȁ�K�W{��M�����}3�˝_���K��O�I��	6��'�H[C���۩���n��E�V%-fYD�C�@<Z��q����X):FBD�Ƨ])�7��:U�͝��d���Ym�'�eOj^K���E����+��~#����P�����a�����I��7&��(�實)Br�B/��U�@��'A�
�l	����,�N�:^��v�`��� W)uGz���|f�ߢ�[�S3n�Ƶ�j(�p^ύ���<&��!�HG&�Z@�&9�˹����.����s�_�q3�/mŠى7�Ѯ�ZQ�}�i:�4�G)q
��V��x��F��	
�y&������K���y�~���ɹ�v��>�����_]W'Lx$[]P�sځp�G�bDq����i8�[��k8}���o�,���9=�H����LB�����Zߡ�=���ŚF8Z2��Kn8J�H��vrn&�����@�D�,��JԤ�|/L�VEx�ϛ�V�J�X3�}��K����ma��j�A<+�fq9͆�^,�a��$�tw��w�����p�?N�%h\��q��k�.,�?���ԣT��� 6M հ4fY�e�r���w=�	o��E�Z�Щ��N�}���r���V�js�Xٱ�w��vƥ�v��wx��`�^i΂��[����A�)���wĈ ���a}�
���w�ⅱ�[k�,۸�uQh}S�M��f'��+I]M�7Cy�q.�4�eܴ
+(�(�<�Υ8�c�ɺl��7���;W���g_��ԝH�j�-=Ʒ���y�S�{��[;Ch!O.A�i��>Ăx��b���{:9��P�-�Af/�0n�s�rd4�hnc�z^q�J	*�T��͜s�<Ԕ�W,�{W7���ת|�!�%�4��vgȊ-:^���?���^p;Z��#W���׫Z)̛#x�����|]�{-(&�o8v(���r6��6M�V��?[�;�라������z^ �"�8I-�-���d�%���% �}@��p0h,Ɏ�]}C�l~���ThSA!qy�aֶ��ے_�
rS��#Ƒ9�ݑ�X2ᓢ��+%����Y�o,�;P`#�"��cӖ �(h��/1!2����kJھ-�5q�>�(�/���<Hs��R��pW�,b�v;Cb�yk��d�ڒ7Z^�PmG��Nƽ����߄T;��֋���>*ET�[	��?.;�J����7RWS�y:���/�k�^w�%�����';"2;�u�U�iea�\8 ����=^���K���u/��e�2G,d�$ �6JUܒJ5:
��_s
5��$ĥ&� 1��D/w�i��$����*��Ǆ�"��㏔"��q��Ϧk/Zȭ�������Z ���{�C�7����l0��V%�>� �h �[�#�+��]qaERQ׭�~��jD@�V�DTy�XւZ[����ϼ�5&}�A��'Xx$=�q�/@��t~�Qa1�
�u�Sr�	���i��f��N�}G��2��1u��R�#���_��"�o�q�A�3��ޏ�?z� t�H���̎���A�g;��z�����R̂2_��sA�}̅~��I�&8�Ǆ����ͩA��~�e��E/�Dck�y�ܣ=.`�t�xX$׷��K�4�./����.�d�t����[�-h��`�|˔̶���c�[�R����1|JQ���NfƯ���z[E���&Fl˨��"mG��Tq	ލ�KS<_�,��v�=��`��]6����莝P+�R�ˏ�Jkș��:{e��[�~MB�N�"/@#�T�m���j�#R��F����Z��63�$n���ɳ��䪘��~�{hPOq��TK��+�'&�|���h���;�ӅXIWV�b4�l�����H�C
�r�l�)e7�
bQ�>���<\YI�ic�Iqɔ��Ä��s9�P�$4ePҨ{Qa���?���lK����Ģ���{E�>��!mK���D�~U~���>^3|ڹ@��~�����Q}��Nf���0�C�����0�ˑ������u�K�8�I��YȂɀ�L���H9�����@�I5����.�z\�T'��(��қ�,-:��A��d02�a���+�st�G��X�0��3�S�ۢհ)�!R罏Yv�x:�����$�����D����x�U<�ʭ�<z��H=�H����|����O��˽�R�/��Q��*�b Z)�4�oF������Dph�L��*?�bYQ�Y<d;�lr��㭏B,n��]�������0�N�R+��B/�N9�ޔ�-�gRi�'/-��0ag����F�c�C����ڿP��[�s��(9R qϊَkb���2�hh!&�G�ϣ>���8C�lʦ�9'���=!�(�Lߨ5�<I�ö́�Q��\���H� ��T٠��{sz��/�O<�A�w�"�<�̱Z������VԷ�.F����$\da�~C����iOV��Ev�s9�p�º��IU���*HDTU�� �Y.Y�Y���M��,�`,��ݳ!ӈv������if�i����Ԝ�$��wR�Փ��7�=��+1��ub�V�ۣ+������m+5u��1[�x�2��;s�c���j�IIkIR�"N0S��̦pr0pj҆w��kQ��lo�i�'���-�%a ���%�z�V�ל8s��^n�	�991����pRzv`f0輘a���f�jt��-՛7�m��ң�b/V�M�寎���L��ꏁ��Qa�u��[�����2�"��C2�nq�$���/���l*_Crv�����p�6��u��L���g�k�Ĭ�F�`�����������c�P���y�(���?1�\0t�"|�HC��*u��A��`J'ǉ=��Sblu�V*tA78��o���;&�mEu����~��6��z�=n��w�O�2���A�a�6�UK\����aeE#]� �R��:�߬�qsy�#BEҏ�in�ǅ��)H^���'�P���2�}#�$n
�Z�β��u3!�A�`/)��^)G0��&���9���[}���4
�C|�W�/���;\�ݧ�AP���g��n��� ?��i���"-�?������ ;Fw������R�&7�q��O)��(Q����k�l#֫�.��ه��	���Ɨ��������	�Mz��Pﾁ�J	Us�~��9V H�	�"�b<Q{�^�>�}�*�!��d7h�g˙��B�-7r�8���]Y;Ŗ5$	;N��  s���� �x�y�˟�$ �U�S���-�T�e��2}hnI3;��q��Vn��!��vP5�1d��G^_`��u�����k�U�g��/�_YMN���l���
r2"�$�x�í\r��-}9	�@wlϛO�+V��p�7j�;$yyH��i�@�'��P�,e�|�N��1�TI��`�F`
$/o��C8��Ҷ�_���$���*����kwR�T��F��}.oB�l!:�o���q[�[�}3ҵ�9@0���`�+yh	�Y$s����嚭��m��ch�r�m��9s���|���k��0��[H����rW�n���5=]I�����+�ULo�� Ѯ���	��p�/��G7<I�}-��j��Y�Ic5���c�X1��'r����=C��7�2.��g8a���Pe�{?�a�<]�wW9�����ʆ|��P2Bڦ�137��'�0:�����L`�q[��AJ����8���x����W;�&:*����P�LCj��&�����|��c�X�%>p�)a�,.�N�bD����;�y	��k��	q7ǫ�9zC7d���U*wc�֗�r&"A��,l*��¯X�ZD|J]`�LB�T_�d��Sڝj���e�b_��Еc󱞈:-�-�5y�[G&fB�"���U�^!�,��pI+,I�5�tlv�)�~�/�e���6Q�{�h�Y`,�qrI����,?���#r�����j����Ii�x�N�X�@�ȸG;i|���^���Q�$!T
�8#z
[ןU��fG�2_�.Ki��s_�C�n��y��}#���b��f'&@�ѣ��[#��E1��3��A�`�2�='��t���D]��2�`���Z��&t��_����)s痴�[H�O ��@�Fw�Jk$Ѝ����Ϣ�`KҙŹ����^%ιV�U�-�uS|j�p��2[�<�zh&=_�Sߊ�p�8�k��B�����.�s�a~��h,
��XP\���? ��z	}��>�,?0�z�T�;My�t���h�Q	�n?���cߘ�
cj���	$���u�wX/*��]�:�I��0�DdX����2M���}��1��lXK�i�ň-�<�(�vg��Xt:� h �D޽`�vϧ,��
�E��͚��n��݄�l&�x)ɐq�Qc�\�jiK�@}�p�o$xfٸPI�-"Bo�K���k�\X��7�T/�#��(Y9'?��+<�V��󀝘����nLb���b�V�"��/�ٍ�i1���T~Nz��C�s"h�8;��z]�@joL�L.(a/<U%�G�/�:�eR�
���w/���6������7l:��`���{h��T����-Ҝ^�-�L����)�&7�����(�G�QN��f����yu*�7�Ҿ�fh�d��P��`�kNΜє�g�}��n����;�>7>ܗa#h�_jr�k��^G��kf���"�9�uW�A&� 1��1j�u�w���լ/�.�}��&z5��1�
�K�+��L�ڊ0q�p$���NSO�45�^<���3�5�ǆ�"9�c@�u]��\$}�Fo�(���# ����S��e;�ƃ?E��{X��H��a���-� ���J����c �-T.Aϫ��1�cￍ�t�R�A�4)&3��O�"%4�����
�M���g�p�?$?\�j�ͽ�l��M�Ѱ{d�^�3Yg��<����X���G7�d�$�u|V�BPg������~�g�.Db�J�Q��86<?.
��A�@��ov�����~�'���͘��C�$h�,IQ#��e�[��JJ�G�M�?I���@��C�@R>�R���B�M�_++�:��	�D�VX::0����mY�$Ȝ����Y�+s��orJᖉ��&�,�+A7���4��6I{�����m !��"��U[w�d��k[X�P���Q�ג�\8�$� ����/���L1h�g��0�~0$*m�f顕�l�a2�7}��p<�h�}e�Cf%Z��Hz^W����f�#C7	���y���S��ww��3Bn2 ��=6Y�|̬9b��M� �6{-�nDx�3`��,.�:
�)΋P�>��|>v��0	]:R��1�i>m��ogO�7�ڠ���4��M�T�<��!�:�Tŭl��2�H��)b��iV?��=��Y��N����ܘ��CT�c���" *폱r�D�-�r<���%�R�XE�5�5��WR�TzO�Ҡ?�r�	U���R�q�Jq���\�l6X���{J������%e�w���˷w���<�]q�|]a`g0�E�,��3�
��o�Ì'2혟�	+���8�����]Ŋ�*(�y���C�1r�.w����V�A(��]���z��klT��� X	Y�誘�$/l�'ǭ=r�xzW��/8�t���g��`�B�ߩ�p��Dm�S)� J�Ǉ]�=N�WX`X����Q�\�<|��ߓ�hh�c�XΚ���Z�"�o��Yݰ]C���9ˇg��4�H��e��1�iEњ_�R3tG��f��!�����������f?7Ӷqu�\c*1g�u5����2�Ii����^�����ʫ�7�(�]�`��Gٜ����Ն��8Ϗ��ֳa#�U��/�I�f��"�3����F����q�����ԑ�(��p�Y�H?�o�7c��SP �Kh]|0�P�!H��AȾ�v;�R�*������=�~�]�a̓DnH�,Ȣ��jR9�=>�{/$>��^�U��A`
P�b��X�4��EuG����ʶ	�O]a��$���	t��a��%���H#�C� �Xn��[,��c����C������H���=�ݑ��.%�|#
���ol,pN��Ӌz~xwݬ�$m/MY���S휱��e4SX�l`��g�6:���AG�i�_���o��͖j>�`@m�����L��H��-��:5��/��X�8I�H���$*��	�r�0�j5k]u��bDN!m�S�1������2Hs�c���1� V�v�H9hmvm��0��z�������!��[��	
}˯@��+�}O0a��_ �M�W4�_\��� k�1�9h�5��N{:#?V3�TRJ���-j;C�rn6xy���g�7��.H���;2��d��jm��R�0�ȝ��6�����y;�y}YDҝ��SBQ,5���H@xW
���,쀬7����*�Э������˝ł��H�h�&٣N�������^�����"�(�S�m7x�(JZ��pb1�s�����!�Me���~��a�A�jB��|�w=���xU��z8t\�`���X����$)<n�B�?a�}��q�[N�	�l��^=t�%��֮ҽ{D`x$&q�*��:R����� Nbǿ�)��ޒ��I?�n�*�8Te	�8�IWJ��~�,%O��fa�QX���؁b�Y1��W��*��s'v>�R���1{O�pM[L�|�WJ�rP�Q��V��tŌ57CR!��K|��N �pkL-��(��;b��*ݞ3[�m�b��.Z�� �.ʌ��y�osC�.��@�@����qI5}�SJ"�(�߷��	�Ҩ��ٱ'W��/	��R����[H��T�Ѹ�g��'`�k]�n��N*�����/�����7��=؞5�$X��^�n���+�6�~?�%�r��BAe�YpiEP�H�s�����i�І8j;���c���c81�oa�W͆���� �YAϒW)���a�m�Iw6A�j.�%::3������X[Yj��9�!(ᓇb���1]#�?���v/�]�+�V��T�{ѣ����3b"p��	uqw(�<�B�c��ߚ�I�[�^�y7k8��E��#:��Nv��+eG�$�%ޑ��ƇZc�	js��~�����s�5�~����� �A�[��ۨ��^Ȋޒa���w�Q�L̀�\���9:=����`���wa�P��	��N��.?=,�P -e_������M�"�4��K������2�(!`�����6��5�����9R���)qƴ�S89�y.���8��C4<�0|�mq���:1Vj<-}.�w��M�N|�e�]�����O��v�F��uH���Vb2�ی��6 àaB���9��=���A�蹼&`��K�Z�lނu���@��R���a�ߘ̵��X�;�'J&��q3�x�5pιZz�
v�0�"Q���m�+�}G�v6�q�tC�����ñ�1��6�x�����O/�ZU*�����WO?����0J*�K�h�J$��o��>�@7�o����5�ţ5(V�{e+�s����̼�!-XR� ����Ts#����H('p.��q&�(���X�a:@�>3|�$�@�i��P��!�� ^>9֧M�Ui?��fԈ\gX|�����<����6��l��@���~(&ܕ��*�`�s\@���Mk�������;�����컻���{�g	�jV�RU�����z��tDČ+�漎���6g��Z��rh�t|�����ő��F����-H�����
|����/�~��Ѯ,�ʇ��6����8��ۡ�x˖!�|�_@�!��eܰ��٤���O�^hV�@�z{��Cb�m����P|q����I��Q���me Oc.�cp����v&y��B��k��1�<}����� ��>�|Xm@��"�u��z�_�A
����x	:�h���&��G�;��g�F+[1�Nq^�HlJtsYr�B����ŏM��s&�.����	=�?��9��"�D���h���w�^��F�b��Y��r17�!���Z|[��E."@�����Dj�27����l�PJ@Qb]]�KB����4@���i��K���<��Q��&%���=Oܷ�Pb%�����-ӤGv����K�����^]��:_R�e5�@H��6���"OƬ�J&��j���Ɯ8M�\ծ�4x���&�fU4z�{E��	nq֋[����z��?cP�>)��Q�9m$h���?�'wI4Ө�LbT咿,�;�)������*R��O��>w�]0�-�5�o�QA����Ƀ(��^��BQC���-�	j���C@���9=]��u�)[�Iؿt�,$Pfr�aL��@����sJn����:��P����՗Bt�Vd0!�a֗H���>0WR��~5[����p��Z�ό�A?�U�BT���ڂ,�>���x�_7�]�i�Wh�?��p{NcV��&�@��/J����9�v�\��)�\qm�s��F�+/:�F3ɲ̀���^�������9���+����?�����%��UR��>���e�)�9��͋��z|�� ���\�q9?s>?��|9�cuMh�������0���<*�`�}f�H)�L_�*|iW�'�\�&7�Y��B���BAA4����9�6��V�L�������O��~��^	���������\sYI��4��6��N#���q5��θ��ݜ�r{\�lGl���������v����2�'���"��*���kN{/&SZN�e���~M��n������R�sU%����m�R#/���?z�T��y�6��ycC������
ᙺ�X$�_Dۋh_{��D�U�W&f����;���j/ƞ4�&�c�FQ�����J/�����zV��e؋�_ù��i��c
!����IQc���c���7��������9���O��^ڬJ��P�M�������c�!���=�4�I4��XX��P,��}���t�a�Wѐuj��r��Z\g]TƎ,�D���ӣ(���u�t�ܪb-��>�7i�O� R0����N�$*p��_�@�����x��u�P9�;�g-�	躚j��fk<��m)��!$��k!�ųτ~��ɢ$�3o���`���"�	� ��/����=vǋ�O�F?l�	��i|^�T�[cN�c{[�F����L�Z���h�u�U{�^�daJF��`�.��i�yظۺ�Q>0(��}��ޅ~��G�1��Y�
�x������W�i�H� �[��F�k�m�h>�s�n�5�G�����Rg��NGc�� ^#�T��{A�TOc����D���f�&R�o4�;V�d�\A�Y�c�f��c��w@ p��*_�f�����4<ihSX+��#1����?#C'�=V�������s�8!9��%&H�Q�J�|�O��D�@q8��%+�{��r�'��dF^у���0*�k˚{����%T���"o�O�H %��1D��h�=�G��
e�ڰ�����˷��~h�\��w�!�����Y�B��l�E��8�|̆{��#K�TiBM�� X��t�-mq{G?�d"G�+=��r����9
ft��
�5.{�n�H���曝�I���l���$�"����C��}���ͯ09ۃ8�$�m}���<��g��'���뺫A#pw������/=K�o�>򺾹��0ö�#�4��[�<,���W�|������J��ND.��TI��5x�)( �N��K���h����qj�IY���g�[(�K��}h>,6O�5�x�܃ Q,x3Ô���uBt��ǫ9)b������O��5���5�k�E�Z�S���܏�O�e����Zwt+L	���.u#��82�e��K��ee�9�Vg��ߝ��1�.g��}�E�Z�r
>%a�e7�:�}FxQ�7���k���\^�������\�˟��	1+:+g�5<�1&z0C\��Y�٬��1�q13r#Z.��i�ot�,v�	� ��z�|m�|��=(�����S�Ç��q@�X)�����(�Hw�Pit^:�~�Q�C�}����h	��^�:�p4�HjI�0�vz�pW`��v�e|x�l�~۵�w1�h��I�&�*�B����U�ثC�v����[�s��Y�#m�XlcL�k���`@��)X�llk�#A�|v��Y8�J��	U��M� Q�fS�ם��h�#��<2i'�wɘ����.Z���[ڢ�x� �؅1q|�`���~l���
.I�ۡW��N�'w�*s�h^�?G���hNk�q,S���Z�C�(-b�ŹZ��3��r[��J�ۙ��s�e�Z`�~��ՐRں$��µ�L��/(֥M)}gd��{{C��+�g�p����|��<��D��2/()���<�c�0����2S~���)����9��!�N�S��v<-)���o�ҕQ�P8en	/�a�9�NV�E��'�'�G5 �̀%�G�:@k��X��K�~�qy�́�R��9�!W���(����BRB?!��QY{GI#�.#mqs�8I��#���A�M�ܸ���s�5a��9H����}>��@������;�����#�qP�B�Rq��4�W˼֫�ټ~�͒���vk��j�:�6�iJ�K�Dx���b��3b�:T�_%���
U�i����́��
�E��
��"���Zyrm�.��3��^���8�]��Tys�諠�}l	��-���F�N�@����X�gV��~������+#�d|J�,�����������L6�S9o�=@�S	�P�܆*�d�U�S�n�]������!.Ɨ?�,� �-$l��G!��t (>:An�����"�(�W�ԙȯ� ی�]�o��7T�wg_f��f9M�*�a8��Bԧ�&yv�E��-M_A�|�&������hd<`����)�u,��+��z��4Z���H�Ň11+vz��7�����Wǂ8NA��l��6��
�g�Hh|���B�<��.!625��	Hi��ۉNߵ�w}�͕5���tA�5�=f͇��_��,�.�q������N|���-��C�B��j�K[|^��F�D�ݕ���^�]>�5/B]3V��]��C�-<�\���/`�h4��F^��n~���n�:\�F��(�*~g�O��Xl��ʞ�od���,vF����aSz3@[�E6���_SVȻ�K�h�R��1���R�a��w֬�?>�%�#\ތ��2G{�і,"�� �)E��o�o,؍;����=�1-��2�W��I�,�|���^����>�[�˫Ҳ��Dfac���],�ђ0[���S�}��DgеT塨��~8D���@`��`v��-�1�d����x�ão�wS.J���j()V�<�EP)N�#��w��V����sc��_��a-���ٹ��E�(#�?�����!S�Γp��U�J��W�x~e����s�6BT����ޖOu�.��^	jgwc^���F9,JI��4���ȅs0&�	�ʤj��Xҩ��t}�uHƉ�,��>{�~/hj�;���8�|�/�,k���L�p~vR�~P}�SA3Z���򾹣u�8�~v�Q�?���<	?&Zԍ�d��v��}�s`J����T"�P�[����Dj��H��ft5�i{��������w�o�d|�hԳg�V�eX�ȓ��~�qx�kC�\b� ���TǊ�v�/fV���y"�Fw��p��*��9<��Hc���FT~8�.�=U��i�fQ����x+F���.����Wb,��C;-�|���^�i:{��}�ɯ��\�S'JȪHt�����~-��I`�r��]�dıs�FD`87��:
�sN��}-`g�1���#��ˣ�p#	d���$�%xr;�x���A=x���xq����Nks!:�Ř�-���J`�b@ap�)�6��u�Oo>�$tf��b����w03�O����b"a� z���-�5�q͚�ek2��?��np.q�\�N�
���[JI�����-F�A�Fx�pwO����C����HV��g��L����{�k��-�xW��q�ܵ��T%�z"�~#8����A`!���ğ��t/�l�#�$0{�;��uaw�%:�t��@�M��`�%:Jc�[1�ƕ9������粇�j������[+IЍH� ��Y-�+iK���t2�[�l��l����?A�<���%'g��>���#;ݑ��݄�^}K�鯀_Jl��,ˉt�	S���m��v��r�n2ߑ@V���gZh���<��A�����-��`k�2�U����`����`��x�2�JE�%.X��f��x�#;���M�~��J�(뿾4ٛ������r�P������%u@m�T�:��O��+�p#N�������� إ�I�P���1>�k��!%�E�z� �1�sPQF��1ա��*-�e�{�(� �`��ќ����J�bj�]�s���F>r�� {�w	o�/>��di�~UxI�[��M[D�(ܢ�E�=��
�b���		x�|��UgW�b ��m�~�r��Y�0<�w�(Ifm��A^���=��E}��<�0�uz,If�CR�S�^�=�k��M�)W�t�хY1J�?;���)�Y�輏��n���>�FRK�ch�
CPB@�0����v.zLr�:D��%9�A}�y��R2Wv&r
�Uz�Վ1A]��] ����&�/~��6}̌#��;`D2��#��<�Y�g�Ncz@-�&E{"��ӉmCRy���9S��B����U��=FM+S����m�����Ŕ:w_ �����aW�,�Y��䀹�.F��h���� mD*�;����k���[�츶�",�Ws�h��K�#�� !���@~1M1�����W!�3$D �P&q��H�.`c�����H�4���|n	����{���jDwn���|��6|s=�)��b{���"p���epk���d�~b�_v������T�����w6�#.)ڐ�S^�2t���>	diYu^��&�}�9���~��vm�D�T��. 0&Rع0PQ��]~��E�*��Za�`?�Ie1�{��=�wc�����Q�[�]&2���͜���
{|V�h�O��dk��n�Cj0mgCQ���z�/G���0V����d'�L��Ov�:�N���lC�x `�~����T#z�F��/��{�)[�&9Q#޾���m���0����˵i�_�''�/�W��FGէ��]�f+�S]��j}��9�΍P<�Ѐ��:.�����`HX�| 4
R��sK-��6��
�X�M��SC$=-D~H�@Mo�{G��:�N�T6Bv�|�u?<����z�@����q&Ԅ�eX	﯅FN�aݸC���Ȣ���x���w�ƿ���\H��͠��:'�Q	��<V�����ov+�S������&,ﲲ�eXJ~���ٗ�B���Z,��ͻ��^�.�S�i���$����,%/�A:���Uy|^n���zފ���O�)�t
�L�Cb�؁ϙ�4xX�Ѳ�夈t51M���jV,]� \�^5�{	� ��M��"��T�
J�k@a�N�3��Ƙ��}Dr��%@7䧂�+���/�x?U��"7�)���G�u_:�J��@)�v�`qonL�|V�EW�4��..p�P����cq~ ��Z�L��#�����{���,4۵���@���h�R���Âp�r�HG٬����f�7���S�#v��)�a�>*�tC��[
2 T#^�,�O�tH�"C=���'�W�c�t�O�^���=�%&w+���Ϥ宑�ai��X���C�O�5)�W�w��=�*�X��U�dw��/�oZ�2N ؊��<�3��ѣ|!&�k3&�xB�S>�����w�]���ҹ�Q��\'/O��%Q+��O�e����	A�2m�//�O��B���P�"g@-�����}Bk�1�ong�&�� �4�ug6��qyUJ�t	�TEM�����ng���0���?b�$�����}
U
@o�ъ(!�!��YA̤L�r��B͌l�B�0 �G�68
K�F��2��}�ȯS�H�W�>��9c���k.�9�tp�e�+ߔPx�m���8TT,i;AݛAy��Ij�w��+w�,��̨��?�r��Ǧ���+���ط�7d
BJ�JX~
�"�r0yn��/��~m�ES�q[`m$�I��[�,�R�Aj�� |o�bW�[�V�D�հ�[�r���-��/~K~�����&�T+p���D�'\g��]���T���#t�����U�v���Q�/�1zj.�W��s~�9HA��d���C����R��W;_�c�-Hހ�X��4}�+��7�]�����s�:���Ś�#��ϱ�x��.*ypjdKjf�<�O���KMi�ζ���C�B�ye���m���l�Ē�<<���Y�-fK\�r���*�C-��=[������Ju9#h��*���l/�\
���ĺ���I���G&(�[�ذ�Z]��]�|�d�X�>��o��0�x���:C�x��vg���]���:��W�?Q�����bG�\���#�w���ø�vA�s�(�!�ɮ��Q��;�q
����s�_HI��?y�W,�@����isp��йx�������hU�؀D�gNA��j�G�������F�O&]J���KtV�jC�I�NV��`��4���Wl���:��Ѡ߇*r�E�٘�KG��vn�A�y+��J��,�t#�:2��ֵ����UI��Abo&ƚE�����fI�o�x�E�}�o�Q���w����T,o/�y
�+a�Y�$�N��W��Z>p�m�����
�H�>����/���ÂY ���%�7�=_�4
|~븢޻_KuD��~3O���� �,^�,��5!ᮩ�����I�PM{p����C(8y��ݤL��r��n�Q��ui�@�]	a}I}����R ��t3����J��ݕ����ַ�D�6�Av�9��)B��gs���)p�97�FN_�,늣i�L�l���~"2��'a5�u����_��wh��?4��
N�.Ҏ�I�/��~��4��қZ�>�!*���^��3^����ҝ[h�[��l�>e��-���b�mݐ������k2IE�,P9ݝ���^����L��Q��X��z0�}�P��A��:�ڽA��n�m׆���Ȼ�~��~Ш����[��l�Q��3����X.�������)����e&������$�@�m�[�S�|�c�U��t�O�������.��w�u'`� :���5��)>UN���(w\�[�	�ya���Q�=ʅe��ݽI�cA�0�0���k��;��������P{��㵥j�6�Ʋ*+�:\���ucrO��5����N��~Ǒ�>���>"#�e�T��7/�Y�n�4��D?�[<.��;ב���HP �n�L�qEb2Ks��_�p��ݼui�E���I��v����@�wZ����f�@�q+&N��A�Ɠ1e�N�A��Wk���Q�[ʉ4;q�pI��a������%�P��.�캕I�mC+�o�������='Ae=H)	�d�(RV�N�r���g_�w�W`~e��3�I�a���8E��f�q����~<k"�����k���� d�VE���u`+X��{;�9�����HD��T�����noo#�G�����Ev���C��~)�5�x����%�c�Z��'�+�!�dZS�;��4"�s�|��WM���o����?e��ԪQ���P�s�o3��I����}�]����Xa���!T5R���i"�$�@����%���5
�m�&�P��M<��'(e�{�c��fA���@����nM��О���e��M��W��/�vLR�_�"�ky��c)�©;����C�4��?l�o��R<��~�$�e�3�"���R��P��jJW�F]��.w}�+~�����)=I�h�A���O��ŗ����o�|�q-��-�G�8��j�Y'rt�ls.��OI�1�53���/����ѝ�]���Zɚ��b�%�f<c��Q��X�f��#���_l�KQ���#-��ū>��_㛂�=T�f������ع:��R����	LO�)v+���v	<��ݛ��w��h��3��dI�����)���Ĳ��*�����Mk�)n_��	�g�v;wRBS�5Q�͂���<����\)�gyD����|�Z/Nq� �#�Y���@R�Eމ)&�Y!���f�٭�?��Ն���&H�v���#2dm�4����~w�@2�DD��Y���$D{wCK�m 6R�
��RL#Q�����b#�a[<�a�H�\�w�J^���R��PJ�e1{��`����U�+h�A8��ۭVes�f4�J��o�ǌ�`�	�j���Gb���?��g{��II�!O�`����_�Y1�U�D�ף�m�NVV9JʕU����Ygu�u�g��i��y���h������@5���"{g�`�Q��[x���߄�����R�uH`���O߈�����}�G�X���32nmج/S�O�Ϭ����t���M8�`�R .��e�X6�K�2�L�/)��>��P�Cc���>�+ �O3��3>�Z�}����S�͆�/ݬ�:�'��l��'s ����%� fX��>W}@��b��H֕7tޟs��A��Z��$y=�s���=������b�B0F3|�¬�^G�+K�<�Ö'2S�ʟ��4�:����ϴx���Ƨ���>5�d���-ق��q�:��ɩ�R}�ƒ���P���6D����1y�!�	Yk�j[��^;7�����PB�N|Vr�6ǒ��S[�j��[3B�yK{.֌^:H������n�^:��R����up�p}4p�څ�~��h|JtN>
Y=���Cki�"�E�<�c��O>���l���E5J���6 C�	O���3��!,���|}8o����N�~ώ���O�"�� Ʉ�T�8�E�����[*�_��](�.�{��b~�<�#�ߙ7T�fΘ�(�����q-��+ua^kD>�>c�\Iij���pn;��(�_T%� \!T4Tr�aN=o�aX���^��7Thr�8D�$1若g�Jɠk ;�������FO�)ODk`��j5���p�m��kڌx�R������*<'����!Ҭ�y���l�:���Ý�u�T�loH"�������h�85��b�� ���9��Kd4�u{zPh��{p�#O� 1�9��w�$��1�J��rz��@����y�BIZe�#�g�3�vc���'|Qe�:��1�����"�B��Nlr �$-�,�Qo�CK�_E��iX�EPEK,����Ո�񌀃����'.����A^A�5�G�%}\g�a8��XOb��k�k�0>Cb���!�p��f�TG%�Q���L�Ô2�����3{�E����4��	E�#z0�I�GӤ��[��O��Ą���	Cߜ��ÍQ�̨ɝ���C~R}��ܣ�;ZRʙ_�s����s�Fұ�{
H���7t��Ȥ�������7�����Y�G	�-bn�S��`e������}���u:� T���
�K�w��Dn��"v�٫)g"��X�欌~GO��K�ÍI��x�d����ݩ @̃��Q���'·�f��)Fu>�y�3�������+��׻�l۠�>˔~���Z��$�7*�w�$S~xE���$�@����0�^�����d�g��d/�����*ڡG��P�p�۾�v���M*�GY'W(�o�z�A���S�e�~9l�儹k�c]��'�|\k�%�Jh���ԣ�ΝnFw��Y:Ĩ�Uh�7��$hE��r���(�V���W$�.��Aa��,m��l��)Q�G[N�c���x��#V+�"�"w��x[u>|�vrc����J�_��1 �o谦?~ ɟ�خ��u�B2���(�z���x���!n)�/�R �uYL"s�9U�`ˆ�	��x��j��~��C�,�+�<�l�-;���-�E��M��K��%�����=�,�Q20�WKx�ˠ����������3���،U���?�2î��ܧ���$gw��2�ip�!�aup���Ui_B98g3��������N��nݡ�O����?����������/��k����◙�yS�0O��0{��ۨ�.zt{yx�'����{�^u=��~'s@e��dp�s�Uh�"�lDc!��e�9w���f����`:6�����^- Ǧ������� �D���a�k��K<���U��m2�����¤E.����Q�p�Z�+�m��zh�����I\钏��細/�Է��̬rr�{Qi]�PW�n�^^���i�X�r�H���%��9E��L?�թ��n1 <�ǣ������9�A6Ԝ]��-I`��4/���U.�k�S<��m���ī*��T�������u�@���w!��P�?��&E�!ʾ�/�M�nFg���Ro
9�����	��3�m�)?����BaC5��`p_�Su��K�,H�|�W&��[��Z>�XZ��t���?F�"ڣ��OLM�) � I�A��a��Zb�%A��]l  ��P�~l����:��15�9��{�uj�7
*�����\��xA�z���
�ePD��yFۇ�j��8���c��V%[��{.���MB���B�;���8�d́�xO��~9�Lv���=�Mo�s���~�Eأ<��J'���Ln�b�� ���� |�����Ne��v်N��?Zo�;�`�ĊLDƌ��,��Ȩc����KS���C��hr�g����l�4�fa;|^I�[�u�?�o��j��L+8��{^Rg[�J����U �I	OWff0���s��wL*��E��rWQ��*�C�T&�X>緒��PQY�F0@��?���+����h��?�n��s�)h�~R��+�|AE=������JnTǜ�&C�Z�WyK��'*
��0�(�s��Kk����Z����X�S�m� Wd�ݮ���]�`�/���]���a*Y�C��i��E��C���������u
Æ�m��Q���O�}��n�V�W�y��}��ũg��~�Y\�Y9��{����6Q���B��u[�7��ĹjA_�ϓ��M�&��q��8�jV����9_��!�D#|G�&-�W�zg������t������j�5�	&WU��L��A���ڡ��o� �J�I�Jow��� ���ě�����3���^sV�}Jƅ>!A�Ij: ?�<]��;�{P�����\�ڨ�c��|�I�RѺ~��K%�l�wR����wV:τ�uPA��c��`�7�#�bZV2Ů>�/c�b����Ḉ���A�
"��j��aU�U��Wge��[�)����IK`�L9RN4v<tAh���q95,�q�!�+������3�������� E�~[ޣ�Bl��.�@+jyBʿ@���D�$�q���j�q�#�*�c܄&D{�.���C��i�N�a�0�3	;0���o��s��1��Z��$�Lwb����Z��Ί	�V�"���xD8�.l>�`��U9�,<Z�<�r�Ŋ�'��p☣�P��CQ6��Ρ���������J�Su�`�6`*!��V1�w�MW}����/�R�Ǭ���[{/�S!(�
9Q�aA)�N�g���\1���qj�I����y�e�5.�+�[up(�y���<,.P�锃D�w���������\�cø�e��3K�}^z��YNZ}�`�xe��m5���,�x�l4�wS�U�f����Z�k�$��p�{Cb�Fd���<�"�d��l��=�L��b���/��ܯ��=iE��`��:�}T���R�(�{�])^���xϽ���Y��f<�Z�D6��<P喌;����@�6�rAn�&M"ӄ+��LX�ڃ�����x���������6�����9��A��Q��m��e��7���(&j����I�����H-��"09촁,Ư�4/����˄����~7r�~����-x ��W�^��iÊ���-?r��L-�º��?|~6pgB�(EJՊ/�"�{���D;���y�wN���r��J0���DL��ŧ&Zw*�j��VgU��{���sn��a�Q�D�7Kv�=jz�{L�-��X�?o�J݁}.�ۄ�$F�����V�ML�O�Ee�;�-�!I����|�����Cp��x�����}�s����܊���Ճ���G%�g�As�҈�ܿ���I�A��&W���꿫awj[wg9�:�od-���=	wK���K�*(^��Ic�l֗Q��Ĕ��V���Ѯ{7�{�?S���V��]6��t�琻�\Wd
����R�`�$p�l��]`D�nk�y�0���[2M�/܌o� ���ٚ�c���"7�QK<�m�"�+�@j���Ǹ��]�V��ྦ62w	^e8�%�qDyqB�"�hH�t`c�Ǹa��	?��>#�O�Rm>����K"슪���k�)m�brڎ����.&�7�p��J��'��Z�?1�����0/[6��@�����Y_n��l&і�s�~
ӮF�4F@��KT��Ε�P:��Z{u��t�x��Lsy�@XJ�ye�0�;����x������!�Ѓu���}�TNM:�^�T���dOL��4�gϕ�P�6:Qy��Oh�Zy�JoQ_�(Ӗ����>�պ�B�f�NK�X�������+�b��$�*�*������-t�vki ᬸ/F��ڼ"��Q+g��>&'<^�[~�x�ODy��c�z쇩��sLҏ�H���r�`h��٫�cH�-�8�YZ6F�FX�Mʼ��������/6�]�l�<��p5�5��pSAGk��2�}IX�VNo�H1v�w��v�R�ƽ*��K�ǶI/,Izq{� ���Z^@���\ܼ{�٧�����BS�iLo�3U�}%d�R&�x��C��3���{d�6�xh���g5o�S!����y^U��o�!ʁr��eL¾�0_)hiWu�oN��,��1�yg��zn�;�BcFk��:�f�C�'�IUF�15xp��~��,p��G�)�����֍1�+����)_O�Q���.Щ(���r��[%\���xߵaS�}l�߻*eB�ƕ����>�b(�>Zfio����@���޶
~�%zVS�ݥ���s���'�L݆:D�}��}����b��1��F�'�b����Ѳ�=�%t�}J�i�z"˷9i�-����T�5�.�R�U��"D�&c;���<ǯ���IS�n�-���<���dc�B!N�Ym�mA���>�QK\��tYI��YZ��������58�I�^�Np�LU�-�j�L�g�Zx(�e|�"D�;���\�j�͔�Ī=k�4K�U�?��U�IQK�Ai�����WHz8�쀟���6��ao��"��Er�"J�w~�# F3�����̤�D�6�;=d=�����4������P�d���y;
ԩ�^�x/{�t���!��
��&�_I�˧9��8wC*���;�N�K���m�=��.ʛ��>fG��Lc>p.�@ ��[^HY��˥��;Vܮ��i3�C���哮W<�U��>
�M��Wꟊ#�P
9�)�Z��<x�l�ǆŬ3��9g�����ߤe�j+����wh�|wh��y&�ޖNM��.̡dm+#�DJ����*C*��/ttZ����d��P�o��{�,0�b���2�66GB���tyP}8s*E�R�2�F�T��Ņ$7������E^g��+��5x#���7G��A8Z��v��"��H8�����GS�z�301W��(�����W-�H>h��vKJ��EcT�����y]]�Y^�����glDˉQ.K:��Q���I�
�L���� �"Z�#�$cD��oT�{��䕠�4M�a]����r�ΕQrz�C(���+ьVYPU6f=a8s�T@�`����{q�������[��i.3�!�n���$�L�̵�$l��H�S�?d+V��:��n�!��wp����"����O���+��3�4ˏ������ꘐ�-��K��.�V�8+��H��	�{VН���h:׍��L~�I19s����.)Q��m��d��)�K��%���a�_야�%ܭ��g��w4�v�tdmt�8�񯮹���|�_�]�x*GT�X.�Ku(<�!
����M`����{�^`?���h)���Vm��W_�VZ�V�m8�c��f>@�P��(RW���s�� :r�w:�|M	�&S��6v��~'����i*s�m� H�d�h���z��ᰋB�=�J~�x��ٻv�� IuK�]�� �ju��@�W�C�i>�#5�J9&2�7,���v��1F����o������X���Yv!K�R�OeUa��q���P74�Y�������w_ى�@�0�ŉD��ƂX{���{%��(7F�:��`lAЌt���3��"�N�/a?�B,=�5q�}�nZ@��AZ��!B8�B�`r��1\wD��-���:��%rj 1�oC\�ZG7������ 5
â�dD)�<g��!��*ރ�z�j��F�˔�?���|�+N1����L�5�@B���"j�H^��T�!�t|Ѿ���Y�T���.]Z:�{G�0�ɶ��U=N���d�q���[��[~8ĭ�a��<1r�y��� ���Q���Fu��D�ͦ���v��w��˻������k7�%;����g���~��i��c�Ȯ�0Q�l�� ��t��2��]��s[��Q�0��� ��ڝ�(C��Y�Z�شق��
�#����9��S�<��$z1���)�Jy��*c��/!�%O-��RT=|�:O�E��i�_����_:�M �<��w���2���4�ݛK�mI2���O"�XV���f���O%mB��,K�OG��VvϦ�:�وd{�<^�c�kd��b���K,�~v% ;\�\�jk��%�,N/��Q���)[\S� ]�
��u�6U����S�I�_߬p�dV��UkC)��{�u �6�a$��qSf�)��<Hjp��f�e���_Z���ၛ�O�c ԇx���o��o�ȿq�5�E .�t�@��,TNף&��E���o$�_��H����_>i��-����x�!��\!:h��a:�a��L����&A�1��0SC����@]m��~�t0,�6xej��Q{ƣ���/c���}���DGy�#�������A���.�}?����Z�B�Q`���L�E籂��.��	œԘj��;	��$��ł<�d�80��3�H>i�!j;]��
�6����-�\���t��Q@m�*��E�A��T�Hv����͋�q�p�w l���9�F)^�?��Ftd��<�"�j��a�& �p�v����)���l�ʑ1����U�}7��\dKE&OǗ �a
��l�p+�uז�1'�F���z�#/�"v%b3����A�)j�ͯ'�Y��"z�� �UT_F�n��Vj���Z\Y�N ���i	A��/YN1,�M���>Ťή�gp�F���H�9�Y�3��-�f@V�At��(����X�t��KxrʫT,�a���+c�K�?��x���l M��1���$]f�4_?�M��w�aF���I��^ڿ�+��М�N����'��W֎�U�H+�OYVf���T6�p�*�3I�����w�yn�k9�!zǣ��o���މk=���v%�0<�E��&�t�k'�w�C^["V)��9�f��~G���"9~sFp�����V�I�P���}�, ��J7��y���f i���s>�Vh�K�4f�2�Qᛐvʍ��E �����ju�ɯ� ���~�KP�m�G�Lbk��f��Fg"=pB່�E�P�0�+�͍��j��|c˅"��f0�����J���K�2G�����U���E񇘝i�!˛Xs��0�CgآTG܅I,};��ޱ�����2c��e��ŵ���iǪ���24��R��:V��p���ѩ`猗��K�~�z-pO
eT�ɷ8�t�c�0�W�D��+P�n�����e54fІ}��;>��e1��&���Y�ul�`$V-���*���Ì�b
�ͮ�QB�t�(�4�ݥǻ����p/���C�C{��$�D�P~�|:s`��+���E2�k��`��㼸�J��.��ⴁ\��qR���Uѡx`c�Z��Ζ޸�ҝ'��^�d��?�ܔo��~7�i�F(��)ԡv���~G��3�0�	$�޳���uJ�ҧ�$o��qk���y�fQ���� ��*��~��Ê�m�NQ����r}Wp�LZk5+���&�W�$]Y�X�m�a��#���&o;�Z�z�Ė�Fgq��iA2��U3���:�����IMX0@���~A�j���4W�D����z��ՇQ}U%B����K�/���ʆ��V���,����B����9t7�F��?D����M���q&6֠t
ukK�F]W��1�e�B�ډ)�W!p�ny� )Μx��|o�A�@J�[tQ/���x�9g�M�{�ǥޏ�O�Z|�P�jW��BF�O1�@����������}���>7b�u��|xDz�����e��=:��Q�"m?���\쥵��`b�YE%�I���JH"P��*T�v�rW�Sc�&e\�H!+�k#߅�����\GH+x8�b����}�)b�Wo+J[���h�RǓ�ͬ�+G�"<3Q����9'M�_��O�/lS�d��:�7�����&m��ʾP���S55��b#��>�ؿ�B�@�۹lk��^�C��@x�ڗ�i�2�?��С2~��9�=����S��4)?3B�u38!����%Q�8�a�~g�Xp�����n�{����F�1,6X�5�D�^�Cq�EŻ'Ջb���
�3 ��}jvز��x��NB�����JR/���s0j�/)��1��_��FN���	���:��d _��Plr�5Ǩ�?��țD>ml�|�����fy����3Ї�:�U��p�K����ϐ7cM|�]�De��̢�z����|��;��
���ۣ���T{�$3��	�Sˋ��Q�*l8Q@M����zEo��:�}^?�RpЧ���]� �%�~]#���UV�\�d�^���{0�=*��<���i����!�T���tD__Vۢ��
��Xl-������U[�M�����욀|�~q�u(�NV����mlL��w�v,F���jjd�36�T<�aإ�Ob!���xq���If<d4C=���"�.	����V�X*��窇o:�}X#�����,_!����6J�� ˒�Ǹ�Z�<|l�.L�jh�C����d����öH	6�0���]iK�L���/�奀$���B6*Q�Z��û޼ҙ��}sm�_bl��i�/^�����kO���A�M�_[=qu�,H���1h�-�b�!q���q"�Ϫxm�!Oʄ}�i��fs0�Q�ǒy��l"
�@8B�n0%��U��C�^��ɨ4O�2Wo,R�5��;v[ϙ��Z���N]�l9Cr�ɏg��Ma1_���$����j{�x��=��Bt��ޗ94�e�2-rP������Qu�^qZJ �S����^~D���W�T=�����%�r�FOZ�K�aO����u!����E0��DX9Y��~�B�߱虏� ��I(�h} �}MS*f��$d�v���n�+��!��LʱvHyp�1�g?Q�j����j"�?8|�"SԸ8q��Xh���]�	}����F�q��1�Q���z��z���I�e��'��2�2S���֘���H}o����1/5#$̮G.%�g>Np�q���&�̞��M���Q�Hj֩�fl��Q�7N����:�dxj��W�(M�-�1}��ozcUA�R0�D�B�(4~� >�&�!��.�Jll�P`���Ļ��}(��'�O^�;u���صL�|�&l �e	_���
]kv:T�ބ[�+����[E[>��ڽ�d� :�W�B� ds��&��4���v������D��Qmp��v{Iq3�g�U�C���ً�y�h_���k�KM��F���/Ʈx�O��g�k2J7�މN��"�Cܥl�}��O;VCr�|��|�@N��De����s���6�=�j��k�p:f9P��iή�}G���,L%�����R�)MLJv�	���2=��a������V~T��x���?$�~�.������Ke��p�=���æ��$���G�<_�o�/����kY�&�1�Mfht�����Է"�H-Ⱦ��&'�Hg�����TP�%Ӟ0 ���07Ȕ��V�HO=Mb7�Pǿ#a��y:D�Q�RxӓV�%�{~��lW��m�f'�%�!�ÆE*�P�A0��Pmn�UL�O�, ��v�"O�R���0�1ffihص��ճ�֌��od_o�K�Q��E
�ؐ#m�-w��F�*�
{��T�?N�!��"�&��Z�������K���ʌV]ߔ�$R�_S�/�2�� ��|�F]�v7§�9+��my�J�r�f�G�G��9�"ju�k�!���G;��uςЩ���%���r	�{ǖ���c�#�����[k��w໹V��i]K&4ɸ�usl��aw{��:�f��э+��]��.-�?�Ù>��F��X] �$[�V���:/8F��.�2�- V�����u��� 
Hb�:'�!��|��~*����]�tY����}(Ɲ\>x��4LGZ�5�Wc�& %�����o��c�+	���E<�٪20�{��J���^�6��Ԏ9�{_\4��P�^R܍�~�zT����)��,+����!��}�Z��0r\֧C+ vF.b�m�,2�Y\�
�ܸ�j+�S0\��S�?�13��1��
��ɦU�xԾN鮂�]�YC��&�����#���K��#U6�ʨ���yQ[k"nm�f�SR�h>UxL֬�E�S7(�,��!�b���^�U�0�f^��J�P���T��C����[�l��b�2����H dT�6U��J�wO#A�a�nEu�c�&\��8 U%Wo��,݇JM?�ozGG�������*�>�	�h�#�l���C�����������=v=.��٩\�z�� �.=�>�6.��B��\�N��z��߄9/on��vt��B;�󎺰E�?��4�췂(���=��0�:\ ��|t[�8{����"�?��.�dx; ��������E���Qv��9F����Y������E��0��
������a�)v���;�b(O�Kٕ��]^�_�gm����Դ�Z.���4as�@OE�y��Y%i'�c��uw�7��Qd2���c�=- Q���
��(�m�K�WN<{x�+�t=�wDԐ�����ٻ�kL�M�j�����0����D�ݘ[��Y���]YHC@Lj�U�rn����)(���8��u	Yc�`��îr���u����
8���q'k��A1ȟ	�o��]1�Z�j�kkѺ-A��f�Cnn�Z��
��L�Iܥ1"�qLc��E�Q%J��땷Vqُ �9Gد�Ÿy��-�Y�Rt;���~�8�g0�r��c�DA�XW��'��sgb�d���w��ԡ!�4!ۇ����&�3�5\�!����*$���5�	���e-x� ��q��G�'�n^ڠk��8*4�^��r[{�,�a��$,���Qc�x���<>#MoP��ɣ�*���`�W�Ҙ~UHl��K�Y�ڴ���G\�䏝�e�Q�a����x�	 �C���J�kH9�ƌ������#�����fpp5%aa䢢$_�d\D� �fv�^�	���pj�C��;�j�߄_9?R��;ʮ��5��=������t	�H��*:8�� ��2S'������e�J��Y�F)9G�w���~�O����	�f/�B^�*z~�(n���ߊm~��]��#�G���h���ȁ���H���6��R�#q�(�^���$&�ǋ��I��Kw�,����������	ёW~��.0}����i�%$	�A��0#AP)$�s��V74���Q�ܧ�������-�d�,K' ��#S��G�s�R�A��p�׆���	lQ�$�p�c:��2t��>L�1:�Lˡ:K�8bt^u�o����|�ߨu�h�F��9��z��\�c�˻�L������ЁB2K��v�/}�L�a���f�q�SO�=��V�7��l��ޒ�
�a�2�\G�a���Io~[�!P����v��(���D��;���;�&|����Ic$�/�44��=(ck�۷�B�m�@F�E��D�L$�^�������7֜b���J�!�x-���m���<U��NjӮB`��^8�������v���бr�
"�am}ߖ��L^@0�;%�DնЖr�J�@*��pl�?0?_F��lF�q�-i���T�J���q�D�Y�!4�I��?��v�O;�o1�2 �@�w���ZNN2�q��.kg_�@a�"$)��q��7oJ��bSoh;ۜ���`��~1.���.�|��II�Էn��^2uw���h&�bV�ٕ�"����ߟ�9��-B�OD ���=�}�s��(��>N���=V��.0��e�,�	�����e}�(xʆ�v�lac��+� �J���* �������t�pA�(2��/r������Y!h�n�İ�J~&C��w�V�.T5��N�C^N5���	��l���Y��z�3�K��{	�w T��N�S<uOXJaEu�^ɰ��B�`�2*Ts��3�������S>�1Z�=�p�ؠha�����n�2�ךv�]t��Y :���2��4���I����Q��/#�ı�[�`������h��Xa��=Wa����冷iϡ;���_4��2�p�bi�ȴV���MԳnm�~�^1��
Æ)+��ׅA�5��3�i4j��#�YGV,?�Q����yqi�DD�e����!��]����r�N�'��.R0<��n]�p]ɸ��`5��X�#��,IOz��d��!��l1�|��Y&(�~6������ _R��q�æ�Z�'D����pj��U��8Ʊ�LR^��N�o��ڼ%b:0��`��d�M�i���<�������En|�������v����v�i���j�~���3`�i��A���d8_�<�wc'�Qs[(6�{����:��j\�+�ث�MSΓT��rf:N����;��e=~�xP�R�*?����%/oߧD�Lz��4S�F��A�u+<`Y,3c�~^gwmr��i���3�Y�O�I.m?��0W�ZE�g���MI��2�^��[7δ!͛5������R9��E{� YV�,����(�,�;���բh<��S�F��3�9U����1'�%[i��1(�Erp��@�i����4�֜��r��� QX1�ᜩd}�y��=�J�*��Rj����°��2E�I�h�2|il]Hd�47	�Bж�I_%���ˬ �vm�&��'�*o�����'����F��$m����sj���/J��x�a��T�a<��`[�Fv8y�=r�@s\Q!ߛL�<:uigqp�U��]@�=�cҨK�BR�K�J��`��e*a�rC��5��
�`%*�U�� �����-�n��H���_���4�����U�7鐗�m��tv�z�l�W�mD;���{|��Z������6@d�s64Y�C�l�s�z�%&��H�[?q��C4�sp8��f����vZ���<�P�>����Ր�:b$U�1 �]�O�D��^�k[��(\D��Q���M<���@_Ⱥ����~5F/�S���^*�
}�w���0����]y����}��d�;7���W��> ��vX��]�-xZ�Nͤ#�1?2�Q�a���V�����Rv������q��-�pӒT��׎���7�`�a5��J/�?&���e���`����m�T���-�1������|T��&�W�c�����4�L�ߗأA7�� ok���B�z��;2壍�$!�N(�9|���;���6z1*�sL��M'ފ�c�ٮ���\�>'��J�7�I���=�z=.�"��o�~�Ew;1ib.�/!�-nl����>�� �����?'�h�6J��F�5�E��[��O�>�ˊӰ)%f,���)���y�2o�r;���(9C"d��5�Q��k�ev�"~��׫��I�M��vw�q5�Rf�Ro�\J[n�#��->��h�v�(���_���
�wuw
rxm�G��96ئh��t��8Vd�ڕ�D�|ƈ�\rƻ�1/ޗ8�4���Qh���O����_=Ll��U[J��P��qbUz��)��&�z�y�_�\A?�����|jeW��<7�@��7�7Q�)�ħ�D �<�
���U�\T� an������銪��R�|�A����٭�������M�T�劆r�X���i*��́u��QA�5D�Ó�d�_�
̵/�4Zаq��!���v�~H����d�w;�WO�#E8B�n�o�/��,3�������m}���A��w�HR6lRq��j��g�x~!����h���\ %�{�혘�2xb���)�c�0'���l�K* �Zwo��ʘ2<'��G"aog�tO����)G΄���c#O�*l}<!Xw�-�Wv�q_����97��w��0�uO[cr��$"�i����X1w�h|���صgm�� ͼ�h���9�t�%�0�x+J3>2@�1x�õ�ߊKV���IA{5��>�8C�e�w��Y�Y��!��B�Ȱ�j����j!6V惥���������Q��m��|��c�U� ���0���K�z��P����{��Rw]�fj��{��bn?�s�V�� d<Áq=�=P�oێ�oV�����^"0��."f�N����Ke�T������h�U`8�~�(�y}bA��u���=(���B���>��P�W�6E�����҂Yza��O��Ǹw�@�u�.�.Q9����!���-F�;���Z%3�V1�a�ޕ�	��0$A�I�P�{���FJ�Ώ��$B(�v�w��&����B�VG�um?��6~�����k�/F��ON�Voio�P R��;��rtȀ�LJ!�K/�������jh߰FVB~|�,�-��<#��H?����IwS��i��������-zC9�b�pҐ*׮��aɻ��w4ܝf�v�F&5-�a�������B���e��Uc�l�B~���yF/vb *�<-%�Eg�ꥁ��9C w\.��ߑ��c�1zc�%KSoF_pQSZ�SV�X<*_@�!K�
�Ѥ�.��ٖ�jK��Z����#p��ffG���i����θ>�T�A������e/���z�&a��Y���5�	�k��<��Kr�)��"h�gҢ���1?�Ѿ6��-��v�	P ��6_6)���{>���8�S�D	���ç*A�76'"i�[D�#�J�7��4o����L�g�Zk�g��Z���fH��|&ydY;�IA���d�pͲ����P}g�
w�>�xӿǷ_>�!']��k� ���͆kh6�$QAIEs��IM 2�- �-��Y���J�ə�$M���C��h�Ǩ�������lyYs��>�QXm�j�jCF��nZ�M�/Rυ2�IR��VyCf�����-ma��;���S��.�i�S�0a��5�Ώ��IF3�i�&=�a#�i	�3^����T��3?��*63�t�B���H&!ޖC�̘/KD:5oBi�Ja�$~ǥY':tF�َ�H7R��!�0-��Ԙ����iC�WqqmF�� �i�>tJ��%#e�i�s��:Y�s֢�O��Ǥ&|�T���m3��>
��̪"�2ǘ��y�w�kK�@��f�)��m�ӷ�u�򃑋=�0^~��{C�X�T}�I�=9�X;�8��S�d3���e����a���A��k֓e�s����6?���O���X�q�(�����'�Ǚ�W6_e0��΍w�������s�5V&�+v���ĳE\��2�s(K4ɵ�8���U�s�1���������Ǳ���iE�i��c��'c�����z+0���������[�U�>d��?�(��8o�al�5�F�N��_g���Y��J�q�C	�=�[ҍ��Ҡ ������Jq���-��N��R�x���[[�k���%�����"M��2i��/�㙂���������%����<IY������Ͳ�d�BG��"���9lP���J������2��'�dr3��QM�U��SP��<�K��/_4�������[��v���E$��RA��	=��$��ȩ�A�56�曤���Σ��<l�������P�M��{8���/���9`=�E�{�j�9���Z,���ꝯ�?�93��4T��NF�r;ˣa	�/\NI
fJ`=��ٺ�u }D��uv�i���]�)�I%�P����wQI�: $�W@�{�<O��FZ��Uw�N{��{3̘@��o	�N�Ұv���X��!����,\�Y�r��u�gŏ䘞ҽ%9n�n�r���=_��l�(�Y�Gpzkr���x�|D��V�$��v-rc�q>/,>*R9R�1q�tp+^�16�X��d,��+̠�.�3)z(�gM�
yﹹ)�č��#�3B5ޮ����b�\f�t���X������[?"�O�����j�
���eo`�~�X���ŝ+�A-C��q �2�B�m����vZ	�FI���|�`t�2����?���{�v�ԦX(����.���nQ�L��Pͭ��TޢCk��f�'�l�Lt�NSi�Z�c��V�g�~��Lm�ګAt����>6��U�`	�GW@Dˊ5�ٱ� ŭ�v�����Ѡ��ܭ7R��T�*���&��j��}-���f�q��t/�9Pk�%n�%�;�E�Mb�sz'�{l4g���Yh/�Dp�p�V2&���b��}�؉�94�=n����[ "~�h�k f���p/w��,{-noy�i.URh�8Z������(��M�{�w[��]�����ߣPn�['��y �,J�bZ]�¯LAB� ���3te�Z?���^r���K �R�S�����7kF����8�9y_�	z�J�v�9"�){=�~�OM1�0K{��s�g�/i-�_$��CmA���d�X�vg3R��6d��dP�.ƭ��v�.L�_n�w)��ሓpS�n��W"|ƣ����u"ci�b��õ����S$�O�)�[����
;����P���Ʊ5@��u���5(�d��6���h�=E�i�A7ͩ�-�bt1f9�v�T�64ju���Z�Xe��aUǀ2������Ś�����Cަ?w��\J�&�D4]<^��ӗg�dq�Ѷm�[D���x�{�����Nj8�k|1A`�!o�ԙru����~����6)�bsJ��+��e��0c<��W:{s֫V�F���^%t���p�D@�uI
@�(�=+`�e�ZS��5�(M��`�}��T��-���ϢبH�6H޳�װ#�>݌�J���t�) ����~����d2��)�)�r��̣�xWz3�Ut7I6r�����W�nE��Ir�"��2Zp�������Wx�]	�����m���(Gܩ~�%T�4Gee�3*�F9#��e�y�Q��/r�'}�_��TX�LO緑V�Nd�]Bȥ߹�l<:d��1o�����LĤL�,�Omr�B��0LCUl��Se/�ť9�ү:h����V��*Cp�N�P��'�^F=�:({�0�����q���@�U[��c&�m��:��ߒی^�A�@)���k�v������F���L�A>8�g� ��1h��]��@�9q�;�qi�ȥz�E|�V��^�0->�cJ���>����!.��h�Q+T�e$������F����-��_���{�L��W��Q7uj{��~Lw�>G�� �4��4}���H���䋕��K�2Z�1�/XT�>��: ݚ���ދǉD��Qj�p�)M*d+i(q�c��(�ſG�}����Z��s�ؠ�/�ٚ�/r��Qq�/�D�\N<�J�VX7ߵ��'�z�O8���%Is��963u�(*|�e������?X�n׉��I!�8��3�D�l�㎨�N�9��~��x�	 �.�������ь���9?VXt�.g4�_	8�����mq -�{�$�O�#�"�r� 
ա	
&���嬑�\���5�{@��yU>�T�\x����q����w~�t��m�G��b���z*��=(/�MFk�߽dDZ �u>�yK^ak�{v��wmG%<6��kg^~h�֣���)��/����
�ǘ���%'�S|Xi�����A�5�}	�	�W���bf�k��i���]Y�OcZL5��36�MG��G��9߯��#���{i���U'r��K?ܩ��� F�p&SC���
�f�ίw�-���2'S� �����e�o�{�	���z,��_l):1��`�2q=:H��ǖ��5��-�E"f$7ۛP��-D,ۙP���0���m����SmdE�[)qE{�s�A6z|�$U�X����@ �߂XDx
�T�����x@i�0d�wk���Ucs[k�������\׫���X?�������M��uK��F;2Vdo�;������1���~��]�9f��5$��l��&�����&d1�f�+c�3�j�!�DD?�ׇ�� !�.����)^�
3�4 ��W/U��8��:T`�9W5��tܾn�N�m��P�^��Ǎ������Ƀ�g�|rd()�+ӗ;�ڵlp+�B{ļ�.�X�n��]�E��΍o [�Q,���$Y�'�"��x`v�Mkp�h1\��5 ����EX:�ǝ�e��f;�Uu���ׂh�ɩKn��xǚL�����Y�!�?���-���w���n����V����}��Bvl�P�KSNHN�K��%g.�p�m��������A�iw�7�墽ig�M�_��5�-.�T��l��I�K$%����hj֏��/��L�w�\?i�*����!��4傟��^j���_v��#E�1[̞-2�9�Fߧ�Dx�G,�L�,Q|��v��iW���^ţ�V'r�Y��W�ێ��ٛQ�����u�X�� �6����ּ`���{�\�~?�Z���N�=\)f��C.��K\C��׎^�Ɖ�y�ʴ�(j	ݿ��v�8I��
�R�/S��+NE�Gm���j�j�?F/�c�7���8�������W>���A�3d�����3N����luYK �w.����+.@H��⪴I��$��-�[�A�]�{̐2����A�vN�����A�5?Vc��dg�OΡ�uyɠA���ш����[�t�KS����ӞK�3�m�Ad*ݩ�nT�K�wmfVO��w$�gcݰΠ�p&#p�/}��b]BR�.u����)D$���Ϝ�}��p�8����+	��K�������� �Z�p��V�9��0Q�D��?���c0�u�y�f��dX
����gM`Hyi��:�z�^���ͥ�q\���~����I��8Մ�^8 �{�>*�	R�os!e��v���G3�L����e(���H�xm7���Ҍ�A����+i���$�N"S�q8�_ ��{�A�h��C�kL2+�f���][�4PŔf[�L��{�)kPn�@�e�oH�n�<b��즒PK^�F!�^�pƫ7g�]%�rZ�kL���,l|0}������ aLDro�:��=��r�xsW�Y��`!�H�L^!����z�ET;�GJ%�C��P�Mx�I��a*H}˞�<�y�q>N>���cQ�����}�k��E��D0�tFY��'ך��2�m"�f�36p�r�V����L@�=CY���4��P[->6#�hWƧ�R��WE�2����D�i`ύ�|��>&��7&Agl4T]_1<F{���N�[R�]C�� a�qVq[O��z����������q�Xձ��E J$?�I�W�z�x�&�A�l�\]��`B���yJ�_C�{ϙ�	�93e�N�k��,P�����+}¥�f�:��k�͉�'
��JYVG��8;%tu���C�'Q&�D?��|�`?$�bN~�B���\��u��V< '�,�9>U�!��x�s��{�+�G������y�"��&2ze��JM��K�TѩJC�שr�Pkz�t�d��}O��%����*�m��f���ΟZ���#�2���������^x/����B��r��D8��2r���Hv�~#��4��/;�
M�'��gpL^�4�q�&�md�!�}�ꍏYi;��!#AB�{�����2P�c_�d��!`��l�=q�DU�m�:.I���Qգi/��ˑI+w]Q�pm�~|�r��v��vح�����F�� n��E�����.Cw���稠� �5l��ŵ(P$�����:�W)M@��	�C0�["��m	�e-#f��wF��c�S�f��n���3�+��6E-�����l�(M��k3ch��K���7�I����C���iiJ����{�h.%�L���T@rQ)��c���W���NG*s���KI�6Xǜ�"��ޑj�|�22��R���5��(���qi|q6��._�&�~� �!�f��~��@u�}ov���Ή-ݓ�?��K��j�2��:4�t�)L�oz#�ۛb��0V�c݀8�Y�/����~�z��z�!��@x����|&ba������\L�!p�i>)C��q��ᑶ�N��a�!��!��-{Ã� �Yz;��嘈&fa2�8^d�2c��]�p�7�x�`9��B�q��/g_o�g6k
y�|㫸���U���98}��;�N��QΧ���c������Wۗ�*?�Cv}���>-���U��Jz��\_3(-P��NS/��2o�!|$wi�$J���\�J<h��vu�ɉ�6o��eqi�_x��$�f�K�V�F���K�)�Jx|r�7����!#YN� Z~e�������^�@,o�9MF�:�in�ʂ�J��L�,p1��a&��sJ��®2N����K:����-'��SM��m�@�z�
�����_��y�T�a�M�u	������c�3k3{�]�4�ؘ3&�c��7�U��.0�&����*���a���u\�~\�2R��'��r��u)��+O�;��+t���7��ozi��Yɬ9Yͫ~�H����Ί�59�d-�~A9�b���������#����v~��5����aj�/���X
�˵n)��p�+8�,$-DF�Hx��?�w���ыO��@4!�DM���M���-�3�Z1��mͮ�k�����%B�<Jew���=
r�eWI�n��CI9���@8JI�yh!
o��cJ�^�:l+ކ }Ir �t* {wNZ�Wc�0hwc�(�l����Xp�]���!�Ƌ�?�Omȯ�ђ�9� I��uLT�sL��D������+��cjb"� ��ࠄP�6��xz���L3�'�R;���Nu3���s+F��-HFMc�us��m����en��4�U:�<+��V�5߸H�;�:�ձ%��MKi2��l���r)H���s�נ Oq�ڱ���V�����Ah���礥����*�ρ�
;%�p��<5�ٔ��~�����������h1�R=�[C����O
iϭ�����#��4�������ˇpYn�Ɠlr��,��ӗ���%���-F��%	
�:բ���|�թ��rܼ���+0���]X�	�	����cE�Z�cj�k��Q"+7m��2۲��{z+_����IC�'��`?�Q)3eϴ������O�|1�Tk�]AEbN��a���{�n� ��h���%~*����}���;x.�Ĵ����3�� �܍!�~�eƒ��}����ld��~ǲ��[�gSpw��H޾�r��B]?���XrT�q/430�@�h�_�4I-mCz��v��{<�a��ǋshT��7�Y~�dR:��ɷ!�Y��^>�*�3���^��	2���H�oS�.r���z���|����]�NE�����������t��o&X0o�D���R�z%Т��F?
� (6yՑ��,���`�.n9>�6��@��G�زz����17@%dݑ�L	}�;��GB�s|q��U�RI��)��~��!���������~U3�F�����!�	�#{��v(�}N`�;���qt�qj)Q�P�7�I��Ԕ"�N����ՅJ�š���5�yBb,�X�/��Bvm�=b0N%u������m.�u?�HB��~~�x��:^�%�O�Op�����.�p�{�.�M�9Ԇ�2�v$<6s�s^�Re���~����ѻ�0�ߕ-��|�mn�]�����}�X���TR�@���"]�&:p1�@�81"��ِ].�:X�Л�	Bi��n����x$� �x�7�C}���Hb�;Z���bҵY��T�����Et0{����:�e����l�=��`d-_�;���(����'{�@_�}��s��)*+����?*�ݯ
�j�\u ���q�(f%� ����&����YQ��zF�5X�ʦ��kY�X{F�.I�S���<߱�A�ן��b:�\c�i����4Y
������/� m���38��\
��@��@�z3
dlH����L~���MT���p45��B��5'|��k89��uА�gWj�+�������6�\FK����J=6ڔX8+�we��ffFW*]�q�@TE0����̀�@x-�bN�����Tc		�O����@K��[��w����Éɐ��9������+��)t_��U��m��<ҩg���j�F��12LзTEp�;�=�^\�a�p��4'=x�������Z�&L���.��D��|�LL?? d?k��F�pe�,������<�Ω#F�����3!i�H3��5Fl5�}5^�����&ҽ�����#n����(�
��i*�S���s��E�6/�"�vp�(��1xz�	�����=k�Ƃ�I��RyX'�f�N!�Kdmi��FP�.����A��C˵��Р-|W��.:��.�A���e�$�����³�9
���ڌ��:�}`�1M%�����ly��l$	{���Ï mܙ���&�K(��ŷJ!2,�`{�ç�w�T搶�3^�?��å���rl���TfU-�v�.ew�mH�:�+hh��������cG��5�B�H	F�a5hů��`Z�RN	����9�V�6ŹL�fX ��*U��l��h�0ρT��C����S���������.�[���:	�_��S	��R_�L`�D���٥?�.Η��1N���e'r���& ���S,_�u���MJ
SR��xe�$�fr+�ǫh�gϬNO��-�HK�5���a�f9�a%'�.y���O�b�}$�R�[D��]�Bmֶ�[��4̀��~��E���/�$�Z:�ҖZKw��֌/Α��QK�����nZqm���s� �I2@���� +�ǝ��x�Ԭ �n,7[mF	3����+�W�,�����J�p-����� �#5�%pU�9G��8���T(��R����:0��W=��k]��l�$tEm�Z���y�S.�8j4"��y�K��~�.Y�������^i��L����-�9�)�'�%n;�;$���Ɯux���	�gaU��1�[�T��w7d}�e�FAN3mbV5&��?yа���Wc�8s��1�i��-�ND��!o�@��f�Z]�L�y��S������#���⢪aC�P'�=&�X$��E�[�br"_��x̄F���:�/���F?b�?�1s�֟��e@�{�����h6.����Yf�^��,�:��Y��w)��:1����ɵ����b�9�
�+B� 4;�8�@��!5��������On9�Ga���#P`57�5l�TbUj�A@f�eϪʦ `��9UaTt� 6����ƣ�����c�ݕت��Q��}���j�n���B�Q�*�Gn3"�2��i�1r��L6�8�E�H���OZ��ۚ�=�=��E�O��^�j�0���q���9`��9����sA<@��+���BU�,�H��IЩ���6e�G×}S�C&�^��Q(P�#��!9a|$F�8S �F.�(�)�Ls�f��)��.q�qv:c�Wա!ߙ��j0j\�4��|^;L���Q��jG{���D�r��g<z؁n���)�i�"Yj�����w�JK�BAm��b���7�Z�1�8u=����#��A_t<iY�O�ā�6�����RX�R�O"�c��޼����G����iӔ�-Q��'�'�n�_3<�0��b-�t�R��6�E#�.�3��9����0a�s�K��zm��n�a�%.�����6�]N6�u�9l��k��Y�e	{��Hw�������M���Q!���5�,�|�,#�o��K�
��fr.Nڥ���1�����S�^b�F��Gq��t�X�K�Ѱ\� �Iz���FR�P�����3���ܟ���3�9��T�yH����-n��nPo���#��4��	a5S��B<ҝ����Es�����~
�<�6��1ʜ�7�*A��52$��Vず1����^��d�q$����-�A�ثL�|4��ut&>�b�#������)j��	��= I�NI���1�� �-�{�~��>y�_�e��^�L_O4:[���g��.峦[+Ͱ5jM���]�5d�1�U��?xS���e�8����#��w�m���(��\���뚡���
H]�����$A'W��~[��m���R�;�d���l`5ҷ���F�Vo�G�`����}+7v+5�헁,8���,��n�r��3��q�v�崍�_#��a�TO�1���Vē��
�<�]�T�M�?�(� ){B�1;�9h�*>c���x��!���P���fr��۲�'�$��m��Ya�cC�e��0���X�u�q�<�(���B��k�IJ��-�*!���a����K�I�<���,@�YwQL��� �yg���p4n�k����A4Q�;Y�����&�8�3�+�8�՜������"g��og(~��:�\U���ҩ�����.�s�KPW�����ԛNJ��������~��ϸ��z�<�0�R�3�>��55h-�]*�p�u�9���^r��N�0�b��-(�=��B��u�q�^�3 ���a���~����fc%������O��ڶ� ��Z�XoA�!�������bhJpR%�����㜎�dF"�"�-;�d�b�+�6��֡x���C9QG|-��qW<���)6oꆙ7h�\�/���Plϥ�k_rC3�$�2��8���o\�����L;�F�����u���Υ!�TY�?�#�~���S�.ιwg�ib�K��k�󌣺k�C��lTI:e�n����?�5��h��b�@�ɪ�إo/SD��~U]�D���v�	�[Ep�N�͠O��y�3ӆ����V�y�,���;0�2a��>��*�hצ�mX��4*O�zn1�?=���z��$��?d��9	�e�CR+�F�h<�xW��>�M�7�6�g?����b���%#C��	mݖM:,���'!�锭]�K��L���ms;�	i:ZQdB�,�KɘG�Z
���Кe�X�a�Yr�$/ӧ1>�c8߳?�h��#�gX�tɲcD/,t��ʦ�_b:�o���9R�s��O�����C��:7����x=g0u2��54B�-�>A1?��*ͨ�b�tkLE8b }�@��[��W"���>:�wS���dP�	��m���w�cu�}z	f�r,�*�F�������q�>�C̻���!�m86�^��RsB~�)��Ue��9,��'�M�����%ڬ�>i�}��/�6�Š�x�S�2U���f��C=0<��)̖���_4S�Y<���#XC�����,Lb�`��V&��.�%+�^)r`���+�Tg���AY"6�#}�Ze5,i��!Y"uw.
Eb��_�U���|��y��gE����JL��r��Q�ox�����~� Bc�~?�#����ě
����Ɯ���9&�1L/D��X��# �ԝ�x�d�T����g�(���|�e���!��F�v@in��F�`�Di�99\����^+��}+�{�:���c�w�Cp�Iễ28o���5��)�����Y��n��ё��l��!�w�[D��}:c���j�7]�@��z���r�Y�]/ 3�Ө�P"��#�%l����������\�U�1��g<�%��R��ƞ;a-0��&���~�,��T�)�/��P@a����ϯ��w8,NaY1y�|U�y���s;_2�2z�B���D��]���lzl\����T��D-�XtS�~Ε�sW5��f�y�y�0{���|2R�A�zYWl����빁6�9Uk�\���MƵ��7�8>�y�h6��1���e^�rћ��e8o)�����b��_� ��Rbo_��~��q��\�a�b�{.ކ5���R�:��tx����
=�B��>�F/�
�ҭ��f��u&B!ҥ��^� x���$#q������PM2���TK6�ȱs,ϧ��+՛�T�F�-����-۽P�Z�eo'�� J��r�Um��ۣy�&G�hu4m/�9rʮ�_>�T��C�m;�&T����Ra�Y�3�9� 2�������S��'`��F�{s�;��~HQ��&�.��s�\��II}_�<�k1�2f�"䷂� ���Z䶹=Ʊ��d�`�kW{��J�̔�ʂ�SU�33u��:g���ܵ��>t���G���XL���8jw`�0�����I�Ǡ��B#M����;���.�J<�F#��ꏔV����|�E+�n��h?K����_Q�]����	wQ�*���__єb�帪Y�7_	g�J���|����煒:�H1����OF�̈́�2d�q{����W ��")����1M�x��uD{���ܘu�#�ܣ���Xd���2l�E��P{�b|�=��Ad��v��F����t{'���ώ��~bǈ�=^W�S��;؁A�R��y^�Cʣ���x����N�y�0����I�ػ�W��-'m�i�?�w��v��kR����xA�9��-�9澿�� �p��1��������-	�g���O��_(<�<�lv�����2�"bC�ob}��1TL"�޶5����|�炨c;�$����bP�e���+[*��⿡�8当�<ЃEg�h��z�1�f�i縑o��0�@`������XM�C�Õ�"
��R7��Q��x�-h�����ڱ��õ@j�P8Ѯ��=�.�S�B}u��	c	Zs�^8�R �ۇ:ι� V��]�N5���դ�AN7������}��Q�7��������@������Ҩ03�1�e���������V3`�5�R�Z�El�y��|c3n=W�8���q��צ��j��#�R)����N,��T!��#s����N�!Cx�V�&-ț ��:�Dc�aٝi� \����<��6�A
��l��S����4໶��)C�V<L��Y�k6��ڠ��!���lz�0 /,rQ�l�a)*�[R=ڍI�.O#a���]�?�
9pw�"Y��.Z>�İo��[q�#\������4Wmzh���6��~�{�LQ�X���Ey�ꆙ�Ihr�9�P�u  6)�3���',f���[HL��h�6I�#��&0�ouк�a���u���w���+�[����DE�|\���a� "�iM'���ƠU��a��X��o����^i��4!g�ҁ ��e�鋎�̝*�X('9�/���9��O��6���{q&��Il��+�n�J�7��|Eo|I�����W���w��c������h�,V@oUJik����$2K�@o�',�ѐQN��w�N�e'Y�[�s�M���d���v-���GTщ��_�	{*$��H�o P�#��&90��s�X'�n���٧��p&?��ɏ��M�0bS��K�<��ɠ����$�b]ImpoL�5��l�r�u����P�1$؞���7.�]J���Q �G��i^�]�$|�$��n�/nBE�IR��ˌv�?Y��!3y���r�:��R�o1���Iv�(b�@{��?Q5���x���g�{W̽0]�Y���z�Q��%
�����Ta�oR��8M��l�ՋƪL������>�o�,��&��0Bq���G�\Po��6��aZ�6U�@��ߵ�X4'h�c�W;:o�(v��BA���~�ct �]�/�e�:�-`�ik:~�MK ��i�o�{�̢o�d��;'��	ٜ�}tE%���z	��g�g�@��9�@�cn��^X���~�2�A��z�oY)�#A���A� D��ߓ�h;���J����hE��a�Q'�v�1��`�t�`$(9�:wlN�_K����G�im��zH &hWȉ�Q�ן�D��o�!��$#��p��H�H�^��zQ����ܒ3ѽ>�4	�[�k�� ]V� ��8�Y�V���ɨ8Bz{�:�#�����C�l��.SM�����נU��������0=s��Q?�D?���&�A��H��+���"Jx��K�=z�	Y�+�b�����|������j���p�$Avg4���v%i�i�i�'7ːS/8/$Bp�tv#kx0~G���(�@�eq}�B�+pi땛a$a�aD�2�ty�:���9���s�H�g�CPfp��ͶͰ[Z�|�v�6d���x��kF{�Z0�=11A�����̂JO���߾N%0��_�7�,�v`ۋ�إ�*29����<�|������/����Ψ�B��1!���>�΋�������vxAhOD����4]�1��$�8߂;Ik�sd�G[�PȆ�2e=��9�z��?%�T�[�p��� ��}�d��4�04ߌ�t�O�w���w�>�rZ6�O���;�m� h���7v�kFEx�2���Ϲ� j���Ex4��Y�~�;5��w�Lw\W {W>:��񄹡����V��\�G�1VW��\�rө9M��`h��@f��ay��,$����/�sn�]��hc�����?��2��5���n��\��.����{�|�e`�}�&�x��/�=���'�Qh��@�����r���'e�i>9X�;�e��]�笆�%y��Ԕ H"&����O������3 K�9D�",/we_b�.��w�R�[���Gg�!@�&s��TZ�g��]��E}��E��L5a�$�d�CiG���D	�*�,�#V�,T�<���{������H�=Z{YJ�D�{�t�=s�
�i�D���Cٸ(�6�2�b���������|�5�[�v݁>}�^1�Y
�:_�"Wc�V��x�1sߓ���F��U�5�'cS��/c���g�c�`��~�	���iE�8���*�w���J�)O���Y��Y~�6�]�kªc��즷��筊6���,B�"���j��[�CБ@G��r�q�f�K��+�Ӱ��|6�_P�ޱY)����O�:�pV��)nka�f�p�ۙ��q�ȫS##����~��V1_��p���*>�`����^�uj��U/M���qi�CW�����T���H��9Ѡjt;F�N��n�Bli�y�A.��Q��6cm�GbA��Y@A�7�����L88�6L���$=��g�W�PBcG�{;����ռɝ��o4�ѩoq����1�+���.���j�������3R��R�}R� j	"�6�SE�T�+������*���^�q1��/�Z�X���=XN\A4
�=76���~k�A�1�)��_ut	=�c�� �uxhFD�����b�΂s�+C3s�L�!q�ߪ��5�ܣw�7�Y2j!WI���R�F�G�_���B���:��\��Y����xп��$}g52�EZ�}�e)�E,�hF��K��8!_}�U ا�s^�uZ��MmB��m��@�J
�Utc�� i�z^�ATN��u�)9-���\���Ӯ9�q�E��&��8Ȇ����P��$l���qz�l���(�x·���	�dFWd7�z��OaY](rV�֠)�߿D/c`��Hê�d{��!�Y}�u3���w���q^���~n\N�|ަ�3 v�&�7j�cc���ۣ��܉��hf)�a8s&��;ƭ�������+`A~�U��U� ���Du��� OǛ~�*ҝ�ֆ���k��[ x2�X��9�ڐ��/��.�_B���ܘ���S���
��9��'+�j��޸̎������R=�>�}�˼zWNW$Vh���_X��Ж?˽��'��5;q������/�D��8�X��(�R ��=rv�P������s{)�����^��z+�	`vv_;(�Ȳ�m�1։���ػ �����BF����IJ����"���U� �q�K�Q�&���� >5��H�yj����$�,��&ZB__�5��kD��p8<
(\8�0���87A0U�u'�G�>Fe��AH5�DSi7؏i9���y��w��y\�J7�'�_�%q�"�_�Qٟ��n��Q ����V��*w/Ӎ{f�7ܖ��G`���W�JW��e*�=���ԜنΏ�+�p_Q���Y2/�۞���}B|�Č�FFj�kj���l�c� Y�������� �G%����߮�f#,wJ.b���AކB�}��f[#��zlY�x���~G��bҰ�AB:�CM6=�w�IN�k����l�ދ�m�A���ђ$+�I�%-Cg�I�ҫ�Q��t�R�9iY�r#����CTf�~�:�ib��?ցK�<���K�	Sm����8|W��r�XfL���S��,���Ņ�5��HM?�:G�F*�:p{݈'<��4A�p� -O��S�6��t10��;V��|�b����!/���M��"�L��a|�*Z�'���AB�H��+���	�2�{,Hzr�4���G�c��G�o䍞�~L!�{�C��"�e�� ��ze�xĐ��n��IA�x��{3�y��%C^��-�h����'�.n W�,�9�)G��9�{��H����n�Q�BA|�dD*��ߗ�x`�?݈��{U���nJ����ۗ��j�-#�M��2&j�����y���FDM���^�:�@-�v�}�y�Q={��`Wvx_��� �$�>h!���U>~�H��#2�}Pˊ}��ۑ�M�`4<*�XC_�#���Ǖ�	_��΍�_NX�狳���X�K����D����"Ο��`�]V%t����`p�����(�|u9u��n$�,���kh�=��b�g��i_|pR6}����8�k=ZkZ��ށk�1E���ܫ`F�6������?�AJ#�O������	9
.�o�~�������~K�2�D�l�S�l��#���Z���।�{�pe� |���ݼ��S*���b�1�VwLG�*p�4��)N6k���&�{AΆ�~�T�w/�Q��k1�'�>���4{�y�7;?+˅B�ͯ��!���^�Ґ�Sv�0H���j;�{$�f�ۂ-R��A�%6��	�}ַ���@�l��]��;�®�C�gpZ��f&=��X�6��I��N݅��	����N��IՄ�݈�{/�Ԁ8�O��`;�d0K��!�y��y�	����������:�]��~�3Z��*M���8_�c9��mj�D{^gf����["��N�K���X]�?픳�	�O�D$#��CU&��~�%C�4�1�E[��� H�z2#�"��:Y?���,�糌h}�0��/�-e���ɓ8ֹ�!²�W2�G?k�������r�vD��
@���r�/�S�����-�����b�)�$gI�;B׌.=��zZ�	�jH¶�q�dk�Sh}o٦b}DN��
87*=Q��iR�n����J2!'Y�2a��24����9��@��'�]���^���'���O�L�
�ؐn=āJ��,��m��R���*�d������b`i��o��,�����X��G-&Ѣ�].H����Ȍ'�Uęg��q>��a����S�����k}�/�5�4q����2b�}���S�M:qԪ�L�=r�`���y��Z������=ѵ���c��������<�x�R��������m>���rc�93�)p���!S�^B�H⃲�G,�i��x)���]�wO'���������9-T�Z�Ch�6��A�H��C�"u��+�Bdr̫�8�9y����V�e0��N�z�A�]d��ԑ<rl��5���v�_̕��me@?�� �"#�^�	Si����R���+*m�I����W�2f�c�Q�]���O�ǻ�o [�L�V�:�g
�l�����"]����LN	���!��î��Z�7CA@����i�Zh�����w�0�Ў2'_�	�32��9-����M��Q����u�`�Op����Q�t���i�A�3���c�B�>�	�*�i֪�F->gō�5���Y�Ы�;��Lt,s���V�m�6�TC����I?����8tt�\�Jvy�0�?�7���r
��X��t/�����x��V�^H�3KM����!/4�������ૼ�	�;z���FHo����3 �l����ʧx������?4���n�F���Y�o�6�}�c�8�!غ�jց��+���E��iƑ8�
����ФÝ�K$����Q��\�[�������5a~�}��;��LE}gg�@�!��hv<��D��~V0����*�������k�rR��YRl���Y�4*�����CD��}D:E\:��U*3�����h`NO43YI��yd��+�ʒXC���L�[c3*q+M��Z/u��K��RX\U��!]S0Y��D�.+[O+}،��Ҿ}~a���*�l-�\�M2�]����9a޻*2�~۶s�Ć�6�p�b�����e�x��᝜��܇�JYޛ]{S���nG�\ur7K�8��,G�i��@ӈe.[���VL��$���
y7�.Fg�If$=&$��D��k6�]��e������g�QO�W�-���[=F#y͝E�nvVہ����n�K����j�#����B^��^Z?�ϯg��4	�sRa���<�(�$R�|.�y�'��l�x���y�D��A"�ϭ��a8:f�p�x�D^�;�Z�����ٙ�f=����5&� ǭ�0%��ӵ����b~�MG�P?jW\^$J�J浃09uT��}�Ȏ�Άt�չ~�'�C���㉢� �*���1�<.��2��U@l2�jË��L�{2Z�i?��G�uXZ��V/��\��6�e��Z?�碘�{��G}��,��U�0U��������h�ڊ�����?���wm�g'��l}�������#��ǎe ����˰;���L���7�O-q�N��\6�;O�$DN#��/vN��l�Ȱ�Tf"��z؁�)a�����[/��j�(��d�
�'Ū���1�!��؍����oQ��<�(��&��7T�����Mf]�	U�FTB��$��% x^@9P�??)ǌ.�(�V�� /�_͡퐎�^)wD!~�S�(�&�,ù]K����!7�)* S�{���������O�De��4����u2�z�x�׎���=�P\���\�&*�ۮe�qŲ��=2�#;�|������W�>���M�`�}«>ߛ#2�jJm��,�5l���p�M$�F@E�m���\���#�+�|�s98���L��%���N�M���P���s���r,-��㾵�P��m����Y�}v�>�[񆴑�xe]/5rod3t�I���DeYy(�Y�7�F?^ d���N{M��۳}�a��!!a�JD@W�����"{3����N� LvPDf�$�t��\C��)��ܲ�?xn�fl������$��4��l�04?��$���e�����?7R	q1���(mu�؄�}��z��q�O66�$�����
��r�c��?ե�w7.
B�~��i����� ���JZ�	�_�d8D`b�Z{�;���ה��z�ǫ��
��/���w�}sڵ���e�M����o�C���8�P� �1�ҵ�G��]'2���3�{|*�Ip��t���TB'����K�Bǟ��fO�O�ҍB�g�r~3���VȔ�ߨ���߸�8mD5�n�PQ��O��"m/Ϯ{����v�1��9��n�2�͒
w�☖��!����t��,�6�߼�!�0bR[��kQ�m�W��_7��L��b��Z$�~��}��Ln�O�j$2�Bb�UI��o
�ڥ��l�Ė\ΰ��D�Dë~��YAZ�zw)�Zr8�3��q�O8�`/��K��^0y�YY������.��Yd���rk�<PaQ	� '/%y����~0%Mx: Ϭ�?��Tv��ˀ#�[Z�`G�t�&uWiO\�sg�Ġ�z	�TJ�4�O�H��fK���y�p��}#�h̙��H9E��%���]��]<R�%\�J��l��3�%�Mwif�<A��d{ɧs�\%�x���Ų��6�W]�B�(�� �Co/�������!�� ��E�B�����gݨ��RVb��Dk��~OMS�����l�=
h�[��aΈ�D���5�镥�%���;V��/�ɂQ��W��8�o;i�I�tR��g��qY���R��ip^d@��� 1�H?D@զCiA�T���Y�l��,�߽�Y��үB��u������������܍���a���|�+� `��r�M)\�f��6�\�P��!
fzd� �ɇ��V=@!I�{dݥ�?h�P� LL5�3]k���"�,9�//�;��I�E�T%=r�����I�4>��Q�G�r,_��6��snTu
�G�<E����pϲ����|�:!}��6�@��2U�>̘	�h�8D�C(��#�$*�e��Ҵ0�W ���Y����M�m<\S�	K��ZR�$2�VW�+�0wB���G��l�������n�y��G�#�>��^<�}�Nt�b3�C��oԭ�5e[���S��6q$�9����o�vΜPHG�]��0���,�mm	y�ި�3�њO��UR�ᢟ��[�`b����������2��ނ�{%�ꖩ"������f�^q,h���E�����KD�%��ޢ_$;�ͻj���b��y�#E��wD�}Y?I�=�s��ܻ8�葇�\��%a��5���I���SU�����(�/�F�xW���������A��Վ]I_plU�Z�1*>�Jg)��T�<�rs͢l�3���|8�����]�sX����pr���+߯Cu
����o|�g�!��+��O,Z况���/�؛��E|������ܥ�3G
��r�ў6�W�eˤ�4G!�ĵu����~ �Emo���Y�ы@�8�Vz�r��6.�0�IOf��$WI$���[%�_5ƽ�T�8*���H��_�_ND`;�� R���B��~W��cC4��~�гpF��I>�U�H%N?���+�x�jsb��A��|Ϊ�O.���������:�KP�Խ҇P���,���[�$�`�}?��//ӕ��-���NK�Z�eJ޼w�/M�j�v��\�#$�A(k���=�OOÏ$#�ԲIN��2f��q���p�u�la^9$˺��C�O�somȺg�(�_���k�L{1[	E��k�<�'��l]u��k��\j/�)к��rX�E?����M�a�Nm�7e`_���]+�&�"q�BE�*�^����H53�S{1fB��C�-�n��`�ϼ��\0�
;8����j�bҤ��Om�jp���TZ0oY-�\�n$����/��G���T��3�C`~��������/� 2�[�G~�1{\�B.FN� @�"�Cڅ^�E1��ρMu�C^3W,#��>��}7}_x�,f��ߎssg%�B��g�s���b���~�i7]T}��B{G!=֦�9���gЀ��뛍�z�L�)�t �ܙg��\Sc~�;M�OFm8?�X�J�^��?�i��H��q���׻��3���� �C"��7��K�|>��D���)3X�p��R�����j��lf��'U��,���9Q�mMq�T���_�� ��ܳj�?Ol<�ƪ<�3W��3(��*�6�ܙ{�
��"�FKK�c�4���B�u�
�%t$�ѕ��Fd!UM��r���`��^��]
�Xg��sp��R%ɡ�h�ι.�m����eW�A�>S� ]cv�ѕ�c���M;�eH�͠�S	�Bb�ӷ�P *��VbeP�Ge`%8m��K�� O5����ɟ߲ʏǠ���O��Rg�����O��@6�n�f}�-s�y��8��[��~:b����'+����M�;���+m����8�,K�T��L�OCV��H\X�ܤMm���ҩ�����P�Π�(3�c��{^��S"w�C�l��eL{�6]e��!���|  ���?��	����v7>ڊ��?BT�����C]���b�57�k��?�:�o��VS���B������/������$Sت����<����)a)���� ܞG��X7�y��$\�⨰�?�}�Eʷ��\��Ң�v8���U�I�D"�D���ExLqe�o��=|���q()��W��{���e�CB��)>Z4�'�'=�n�	�k�?WA)F��H�<I���C.�ܠFO�)��g��G�$Uɐe�����mǰ�8y�+s�΂��8l*y)����i
�fb�b�]R����=��Q�J>�!nm�/8������TIU���j*t�['�N��CtDx�6�f(Z��N~���[h��6p�#=T��
�5���Ȟ2F��[x#C�1�"첓(g2��>�%�����Nٻ����Q.�Z��B5+�0:G7N"Vs¹�OڮF�ǜ��=ɮ��;���rͶ9e��е���hW��݆<#ύ�`k��&��R���n��jD]�6�aau�������7:b��o6̝)P\$��m翛�7��e!�����v���MI��-:9��rG)���j�V|r�+�ĖDD�Ȼ���F����|@���an��nd�",��P��u�w< ����Ka�tI�r�ƣ@���G�21��S��[p$��(xMjҜ>��Xr@���Nn�w+]��~Y�Ӷɥ!���o��m�������]�^XM�2N�����Rl?���2��K��F������M��!��p�}�`��lN��x�Ti�t�����/�\ ��.}���nS�����{8q�aq�(�OQ�v+_��N���kQ�p���N£�v텹�B���Ň�d�)�r�� �wk�5�`��>2����)�x1_3Κ��(E#���T�
S=ڨL/jUqd|8 ��=�:%�׻d��F�[�w��%
e���%�U�A`N��`�Gs�+�tm��`Է��E�p���(���HQ��<�͙0�k�*�j�Z�{)G�j���#D��`�L�l��%_.�-�X��(�^��b*L�}�&���f_�עF���4�q�b�/�V��8�e$u��C�$v��1*�tnN�H��m�@k�;8�7~c�+CK�FU�"+�2ݿr�w$o[KM��f��.S��f:��1<�9�3r�D��Z��-4,���c�G�9io�v����xo�l�{��|�\���E�u������<����o(�y�|"}�_e[�h��u�3���Γ��,�3���ַK�=xsq����)�%Fƅ �o��vRY�0���hm����v~�R��e�դg��C��/m$\UY�J �u�=t�
� uŰbi�A����g�ޠ.5���t��D�Q��72-&-���x�5�����{٣��M���=�◳g��*J,�dL_��$�`�Y7�u�*��ė�<Z�ưB�Kv�ʸMˁ�ɜڭp�棗�R�P�P_�y{m�*'�������p���,���Hg�g熐�}��eK]��_�������(�P��I��dq�`͹AP�[��UXg��흡:`�R�,�Z���I�(c��&���"Z��d*�9=#�N���G�z9�n^j�rL,Xl��Nؐ ��)�`���e`Fv���T3�q�]�G�Uӭ%������w�K���M����Q�T!Gt0�(7;�&q��S�H�>�2�_F��E���$ze�X��C�32˙�f;�)�s^otG+����+y��֥��O��E����l�!��7	]Z4�7�����k>k�:������Ԧ��A�Fׯ�<���Klƿ�<�:�r1�࿟(��m��w�#�~���%��x���J�Ĉ��FQQ?S/�Gtډm��}R��bt�\[�������R�5�<c�Uu�r�)zF�ޝ��hLYP�P���C��]n%I܀�\�n�\(���{��Q�S�2z�cS��.���~��88Mj3���gm�T�P�\��[D��3/ZW�j��=�=��c�m���-ݫ�)��I����5���é�v�ȿI-��(2��(t�(�O(��G�IU���D �W�XC-��R@�
K���έ�E��`|������(�B�R�u]��U;)���W�Ы/rf+t�h ��+�o�l�fm�Sv��$�ˀ?.�a��#6(�7S�6�+ˢ֥�.��r��8޵���j �	�^0v�%d�S���*|��T9�Ճ�)�%[���#r׽.?���m@�r�f�@��`Ēn�w�����5���~�Vh�B0Q@�d�5M5�����y��+�b�+��ߋe����D}�G��(��,,������n�������-̎��>h�z$�ߏf� �l��a)���慌Tˌ�-x8��mq���ةx5���j�}TY���qMy�D�}��]&�-�z��_�vB��y��au:RN�Ϸg��nD`�"���U��c��-7m�g �A)�`�x��<��` ��ϐz<��Z�Q�q��tu�IEf�<L������\�Tp���ٜ�x��,���2e���۞��/Z�;�����I��O?������$�P�dN)�ĝ�,�E7�������FSO�f k��J �?�f���F4܎��G��?T���|c�x\�dL1�+ E4�pN�:0�fm�F� swN�˓r���zB���l��@T**�q�b�F�˲�����Z� Z��#_�� 4F�k֕��26�zP���>B���ѼpK��>�.��*nyI R.��_�N좜�����E[�,&��1YOL!�9��[��W�����u��B��s�{G��H���|��!�H'"=�V�v�
kɩd ��T��-oR����J�-�J�;VȲt���	�y֑��QEw&�B�g�:���5�4hN
�w�o���k0BM�ԁ� ��2?wH�U�)���D���v�	S�K�i+2n���E)�n��|���P2��h	��S��`�+oŢ���f��h�Q$�Z���A�|��^�v�t���p���R^a��� ��~˟���ۅ��1�e���2}�P�[��'	���2т|�`��3�K��w�>1jNS-���m3���| �،����L�� ��8�n!o��z�6K�}^|��4kG))���AM�Z�r��+����C�ԃBfi~h��{����LG��������2��rC�d���(/�2����f�F�Ĥ��t;��x�@�3���,թ����R�dV��F/յ��!R>;B]sIS�����Ҷ^���+�֥s˜E�ݫF��DV���t$�D������3 ��y�B�LN�m���fv��P��u�c�y��î��.V�$Q剐�mǫ1�}��N�ף׭m����$�9���v����կ��F$�u�lV�GH����]O�"�V b�R�@�D#[��X�b�|)���Cl�Vo�OԒHU����LÁ��|]ҝ�|�4	�T�e:��N6�G�����E�����v�x�݌Ύ=����L���ݴn�{�l�sۡ��#*K� ���J���H��5�g�?�.�o��h-�I=��g}KVNSJ��*L���e֢tJ!8���h�e~ޥ	�䛵G�&%ѽ�Q�cU`}��Ć��]�|�e�y��e	3-���f�p��z������0a�/�Q�@4���iI���	�|Ͼ�5�I8pF[�N����+�>�M\Ҙ����U��}y�;�8=��^�m�ھ�wD��rsm&�r��5�9Ў7��M�6^��s�f���{��w��N�k���-��N�!����� J K�&��4���u
�uyŭ�0�Fq���2E��h���9�^(
h=焑`���hv��hۙB�A����k������b��zT�}#3�qY2 �u�I� !����/W���e�� �{��|s<rPߠ	�`hLIJ���׽�@G�C��g��� �+
������Њk叞>�	4�郭x��2�;��ی�C�,��39}��wUgI�_��n�Ol�Y�u@�4K��EH���9T���F��3/_ׂА
-�;d�0Z֦��PL�QH,��oE,����W~+K\�.S%j�R����pe���
��۲(�nr�:,���$H��9c�=�w�b��F��Ң>�Hs�����!�X!.���7ǹ�,<�a�B�u��?����8�	a�I�������/�쑢���ee�::-K�
�[&SYmVִ�@k�ӵ�W]�=�f�?��|F%��7%�Ȱ�o��5� NE�dd�\c]`Ѡ?��TO�f@�@����e��58���:��XI�'{�`�F�b�����}so� ��J�/��:(9]�Y��Ǔ�T�-N������@�B7��*;���-4� VX��e�,i��<�{�_�2lĠ��Z�\���D9~}P��k�U���)f�� �Ƀ�d�a��i�I�{iZ^l�x�+��qL�v%ߩDE�Px�F���ܾ�ZĜu?Q�n�Ls�)�|�?v2Ja^���R@c�o�y9���Q�����{��Z=��c茐�D�ͻ�uŉk.�������Մ ���#)a/���ׁv2�zD�3�P��	'x��q���x����a~F�o1�����#�_يt��t�`͝n`�='ԝ�$:� �N]��.�tc{����GY�R�v����@��D�{V��1nwFTc���K?6vw���:�_DX�4��B�.��V�J��dѱ���0�zobC�nîIw�i�^���I�A���~5�����* q��qx��c�[M����>�.&�!�A���>�����WdwQ��{��SuO�<y��u����N��I.�z���Y�|�y���U�$��f��%�lߴ/Q�YIк�Ɇ �l'5J^��A�({�
�#Z{�F���~4���u�;��J00�������)yy������Ӎ]�����!S�I��ǉzNrŴ�ּ�(�R����An���a)&T��P���;�Ch��������I���"e��1���4����TϻI�RD�{��s���@���i���oB��w��k�!��w1�$�KԆH�ʽ�e�b��(�n��A<��w��p0�^u���81C����Q�D3�FT��a���X�$�?%���Jv(f���*mS�����/��RSV\��"����_8�p(%ฒ��]�Sbam(À����aX�r#�ӛ##ӑ���ʢh��^��I��\�ٵM���4$�qd�°���ϩ�ֈgX:R���x�
����[�n�d����k{�y��0�ESC��A�lV�p�0�#L�R.G�(����}lh�A����q����F{�)f��{��-�5@���"l~-k��y�a�u�[G�Pm��q�r6�0QZ�5��QR�&,�`Z��c�C����U����h�ڀ��ʶWMH�Ĉ��e|���:���;3_��4�(����%��5�n �;�_܅$�<zR G�x���LÐ��l�GP
��]� �-�l��{"�괓~�>�y�F]�n#J�9��C4@ h�p�E�"ᾪ�w���B;;�3]�P[�Y�,��j�c� jG����Z���4� T(�j�.�=���|6����Nu�S9��x���dA�	�6��:f�P2�S�eeD�dy�7��Z�@��f�ǋe �T�#�9����bD ����AcaTq삪!�5�҆���R��J�[������O,1�{����6�F�:L%���A��������Z�nPUpeƓ���F�6lk�kv��ҥ�+�Cr��aC�����6}g�����k�֦�@���^*����XJ��vH�"����}�.�[T����K�tP#MW����B2,��u��0�/h"�\��i���ܼ��g^�p;�v�e���qqb�'(�T-ʁ��G� *�~���j"�B�{k��yh�\\?�R������$ptI���[�QɅ~>(�W��"[0�td�,x�8�Z%�ì�W\H?`���$�9nF�(����&=[ m��JϹ;����8����6�_fO ��i���&�����8��A��@v<�V��n��_&+�K:�_�>��qVyMv��Nv`w����r2�(;���P/>t�^H���u,�U���+iY|$~r�W��p��,�R:�)��z����+-���Yf���ܼ6'^ك��{<fŶ,��5�݀k�ӗ'"�\cF1
��/x�e��X���k�X�J�z �:=
�w%%E�=�v`K~���iE���^����./�� {�X��j]��f0'	���M�&��.�T�!IVJov2��E�w����V�g�R⒲!F�V�v�.	E~��`�˲1D�{�>P�������\.Z�M�X?2m=dg�Dm�| ����J�	yD ya�*��F�}��e�*D.�F���������;y��V�xJ�I��i�t���=�?�x���l'#mG���_�i����w��,�3��|��p�@�U>��<Q,O´�uVlż+��FG�Q���;�'�#_^�xf���j��L�\m���cH��=�i.N?k�s����_�!�8_P>!!B�--����آ�ßD�~�6��.�X������NV���z�H���y��E��-c�3W���]F{�$�y~���]�z��5kH[$�p��-��r¶��y�pR��3υ�`3}��y�����Y!0I����T���AZ7�V���\�>#��K��9��0ر��HX[d���o�s'�5�N�X=_��ت1q���\821H50կ��_�(�\��;�3�xT6#�,��X��XXA/�Fx����$�* !e.�C*�ٗ��)�s#��R�m�����!�OC:�����4m��m����),B�ۙg��wX��t�"m�Ӟ���)g�Yr�)�%&y]�UЉkB��D�W�	L��#��܀�`^�+�t2Nx��qOҭ{'Qmzu1��.�#T͌)�"�vtا{0D�)��.�늫У[F�KejJ>8+��yV�ۉ�J�Ph?�� ���v�N	��E̙��p�9$Ec�E� �,�6V�2-�S	���z2y֞����2z�����*�HgC��I�or�?7�̚&�?�S-�Aiw� ��U�v�a���?/��?��]�`���6�!�B�NE��o���})�.�O>[�h�>}O�z�m����a�X�#������ț�P�=+����V�9�bo5=���N2�����b�*��ds8��a�o�*���28;.OƔ���ҋDjBS�s+ďo���I��5�>/={"L92�������y���^R��?>=��n]Sݵ��4<�������$�
}�J��1Rqe� c��yQ4,=UQye�Qq���"�)yF�@�g��zF�_04��X^7o�Y�꺣�>�C;<�e��r{�v5��^��ߐSa�8�D�$��e�LV.G(���Lm�ۻO�?�E�g��X�ҕ��=�p(��ש�h>V��@����qlK'A��o���~"��o軽��h���x�EF #:�(�x�����8���%t�`o� ��ז�(�D��r��䅇 �B\M�8��utt�ٰ��q�Q��{'�W�W���HW�I�;��m�� �|��#�Z��r;s�2���q��)�܀߆x)��U����Y@f:K����:��6-9d�U0�b�" u�"��+�&�2���Vn�>&Ӓd4�~oY' �����w`����`��k6h^�����0H�[�Bl���7��u�}��+M6M�r���͛aZN�#�<?&Ь�Mi;�'u>��<�6�o]dae�s�[���s��Q��vw_�U��8e�Uq�J.���{d?�['@XƛK�Re�*�n@)Z���S��B>��@LO��#�tL<L�O�{��m@h)����/�,Kg増������iiQ�"
�St$u�	(�5��ZD�z�kΈ�����#P_$ך������CE!s�ZJб[�x�0���h������:U��EŊ>�ݛ�&�xw()(C{4��_�u�i@'g��<����w!���,Ǚ6��rm�o�E�����P���k,LZSڿ|�a�Rʩ#���W�=�Z�+�I�hQ��H��g�k$I��Q;��rl5ǋ�b�f����CN���l���6�ph5��3|�cV�l�2{�5�X���;�sCq��V��9K��U���fGO������[5�#����q��ѧ�GfZ����ЀO�[�`�� ��-;�
^4`��4����4j�$(NV�	�΁g�DJ;���A>!�J�{0A����N0o��]�8�ZӒ�w�f� t�2h��+��<~�\��b%Z�B�S��{s��ڿ�5!���̤��2.$-��
I)�ϭƈ�O����:�4�J�f��q�`���!d.�}��!YH�h����f� ���������ދ�z��/o&��W�x')<(Qƞ�2��?o-��:3Q<xJ�Y����њA�Q�MI�A�eDP:Mώ?�*iA����*�z�S+��Z7f6��j���C]k�Ϣ��Ϋ����B���k��l�%����1`��ig.���L�08���jN�N��R'� v�ߔ�w�.�ڐ��ғ�Ӂ�`k�{a���ޭ�eU�iȓ*�8���-���>+��"2y^�C�I��˞��c��t��M��=M�*»�
�ٗ��]��JQZ@��\w�\�+�ĭ�s5#��U���x�yM�nz�m�����S���;���I$YD<d�;0=>��7���Z����	��'�9IqF�8���Vt}U ����D�T����y�l�0�q�ý�e$g�WG�{㤦)L%���(z��vh��(�j�l�����̒6B��h��lK����jY�����7��Y��x�������M�Mp���>��s��@!�LL��!%J*�Td�?vw�5A�gq�T���	_�VfQ��=5��$�Z
�� �CZ�����{.�Kv�S��}~j'��>.5T�7���Xޱv������Q�3�~��;uӋ�j��5s�@9ﮎ;OD#F#�U|��bHw��z�8͐tJ��͗VD*�
d�(ȷ%��#ە�[/���-;8L�#T~�����N	�M�
Ja��5�����U%欘N%���k�UZg�������X�]m��~񇣺����o��X@�!(��Tk����;:�8c!ֈ&|g�Ui�x�+q���޾�;�~��/XU�F�0ԫ����z��LVT�.x��d����mM��W�_�4�_줯�fNw�=�fO]�Q��Pi���<B��B�� ڪ]�[_�uq�;�GM}6hd��q����r�|�dyԝ`��LT���;��	�Ӏ�li��~4P�"-��1�{4^��)R�>>��`uA���s�nFM7�dD*{?q7tB� #��C�<\���j�^k
ڤ������pzp;�`��|��ĸ�M���@�D�DH~��a{�ϯ�i�p0к��/�[�V>9�����d��?��e2��=�=�}D��/�����Tjx��8���o� Y+�z��Ń�WZ��	[��l����[�e���>Ϣ�B�Zّ{�]l�;�瞪MX-^΁$�2�[d�ӥ j8�I-ex��-��2�	lp[�$�����������l�����1��r��C*cy_A
����j�ި�,N��޽�:�������u�p6�<���jp�O8{j*(��zJ��17�������@�F��!��!&���T�e���b�ްJ���U1,\/ �{	���+�^�'@rɴ�S_׹���XpE�k���+/�v��ci���r�VU̽#O�����u�{鋸�[�)� ��A��S�m��?��pN�M�J�{�ի�H��!��&�0=h�JK�!;㥮&�?橆t;,��zDʤ4@�Y�����ߵΫ!/t<�����HLʠ����,�Κ���@Ff�B�PF�x|��Ñɨ��io�i�H'�4 "���g�;ï�+�(�ٌ��[��p��z<	����$�
� � kRWo��o�.�t[̀��av
�Txe����Y��Y���U��ƶ�s)��@tj�"��d��qmZd���r0}0���~t6r�m���K�E�^�	k�1t2��Z���q���Jr�s� ]k@01�%\Js��L���_�c?s��,�06���Aԕn���Y��M����A
^Ev���y���5�[cGc{%�����ٍ��U�fi�ݒ�e�����n�v�b�6����u6`_h|E�M=�%��ڷ���d���0�JF�A
�z�Ɩw�Yw�Z��p7�~�!����7CV�0�~�?h;�-GZ��`�W�uq���W_iK<��Pi=u�m�����Y����(�[�N��0MJ���8O{u(p�C���Π��{kN� .�ې5݃~B�hKL�>[�3�5v���]���� >�Wv�T����H�yc���(F�_�*�ϓ�!���|A�s�B!��br����%c�ƅ��3�bf/��X����8�],��8hd:Ò�NO;���@l;��r�}�f�wQս�����"��Oc�|�#"��H�9���Uo4S+d���;.�4B�y\��
�6i�;+y? ��sb'�.q\f�j-�w�~s�n���E� �Z�ҬD�� eԻ<�э�RעL���p3+r��?/ %M2;��.���s�����s'�~�휕J<�E0��7���Q�Dݧe�-��+���|������t���đ�J�Q�$��s�G<����#D��F�����]od5A�����.7.���+2Ɂ��(��
�S/sA�^�����BZp���Mcb���D�C{w˼�i�{و~��q4��|�(�;�=�jy�kw$�G��	^Iv)��>ã����}w�4�}��inW�a�jt��hW�9�
�w82@Z��ό�c+�i6��*3�OF��p%e�����1�f��g��Y��话"���h��c��<��GB�t\}fh�te"��7��־ٗ����? �����_a��%�A��.���b����T��KT��v
��[�(�㖆NF�-y�$ue���_f�)&jh��+���X]����T�*�=A�ƹY����3hz����b�(�7uه�%׾:x�l�_��ߝy_���ݺ,|2uGۧ?�\8G,leȲ���]#��E¼�,i�ᦺ�>�My`�^~Em����\���A"鰤�/��ϱ���;
K�����|��tn�V��@�#35�����*+?�I�~�"�K���,���!�l!�֥1���ՕU�Y\$5�-�e`�+�&�֜�	�g]�^��!�ES�s�=��>&,�����R�tۀ��ǩ��5h+A�X�h������h��9�Ʒ���ВG8w�Y"��ə�r�n�qn{%Tr�bE4儐 �WP#�i�a
�{��Is�Gmn�R	v)��ݖ��x�̽6}��I�K=��(���$�݊O�%�� �h���]�$�EA ��ZJ�����pT��4�I�doT �ނG�ʦdy�R�|:5����(E���c��^�3�m����W��g�-��"�n|ڝ��Y6��p�k����)2cÓ~?�\~��*>�v�}<6ϸ�[+��b���,,���ر����9�2)��E��SY܌�����K�[�'�v�q�Cw�M�(��$]�3���A�&z�)U7�?Ha�Hm�<�����k�yR�e��ͼڻ�q��]�lK�?���f(S��Wi��3���W��	�U:�����j§?n��o�G�M(!G��-���jiS��Ԅ�8�T�rݱ�h=8����Lꨵ��1;v�C��HS�>�&ӫD�	 8��ѮĚ��R�Gu���Y��P��|%t~�TI��ǋ�*veu8%�7op�s~����Q#S�r�%x�I�����(8�$��=N��hYR����"%�Z�@n.]�YA�3�}��- 61��k3�x�s�{�#�0ݚ�~�\w��9�4�U;�����$�W���ȿ��p�Ja�x|�K����ɦ$r_A��ۂ�׹v=1������V�%J��~���s^�F3! CQ����E��pig���Ԥ���K�>^�(�S[؉1R�0����2>	h&���$$<%�x|9���Gc>�3#
R�ӧ�F�
�N]H/ر�U��j嫖By&�!a�>�/��	c@��R�!�3��b����1����7}uo��I�M�ZNj�du���Y�a��L������+di9�y�	Dk�щtid ��dڋ��V���?>������Ĝ*B� XA��d���e�q4��������a�Ѫ�Б�~�:G�ĉ�zC��ρ�����Ő5�;}�/e�a�
��+o�K��P|��oD�W��c�n�r8#��r*�0��
:������O�iFhp�����S�Q���-E+�>`��L��,�_�=���d{)ɋٞ�,��K�٢�1ǽx��G�����L�E�_��v��A��'��*�F��vzg�)���o �2\���.�!~�$З���m��Eüm���]���qB	@`d�0W).��}rU|xY���k�jTw�����|���!>�������볧/��b�9/n�Y�x��h�; �GRX��ן�\�0O��brU��RT��U�9vQ������\~�T��B�x�� �5~�zcwX?�V)��*̍��B�X�֯��<�2-+�A4�"� ����d�`׃F)Ӎ�ܤ�����f� %6�����õ���?	��Ϙ�(������vv&��Uc���ITܐS��y���ץ_�6Vs��v9|l���[g�����=�k]J�Iz���˻�j���	�I:s��١�8?#��>�e���	�7�hñ��*.L��[9Δf\^u?�o��z�����,��7y$�l�=�������'�B���	�y��>8t/"r���IL:��4n�"K�
E��v
�k�G�1H/@nq��W^���C^o|���/+m�R�ώ��~���7�ocC�m�;/4F��������G����1e��\pF�q�J�ʧp���f� ��j�Ђ � �:h+��a�Od�>�ʼPD딋���=nÚy(Gʭ�����d��V����P�ך�~��M�6b݅�S7DZhX����
z}�]�KYYcG$k���ʤ��β��\�NK8�9���e��*@�vxs���%Jw��>�4��wmG��$��?�w��8cy�Ԝ�P�����'b�T�`�Tq9�@�g+"/>3ր�H��<��վ�V��R�-�<��?a��|<j��uv吭����:����<�����%����]*E��g���8��0i��7yZ����(�*��p`O��T,3��P6đ+sz�<��Y\ǉ��
z-^�U�i<�A�uD�I�\x�k\����$B��A�9MQ��?S����$��ה�b.�����cQd����g�I�H���Y��U8I��D��<����_Eߵg:�5^�l�fh�!�b5�-v7�u���՘j�]�s�+�AI��WoxO)K�R6ea�韂���d݁)�i���?&�`t=4�WY�$�8��]9��G�����o�5J,:�r�*<�������|�l��͠ga����V��:bFx�e=i����_�m����͚u㹟�-�{
��5�B� �]�;*��t*[_��
)iX仏iL�K!b��=���72�r4T�b̚��X��(���lFC!�Txj-�Kخ�[�@m�~,u6�%l�h�^i`{A��}��D�σ9��9��UG#kjPE�-Y��HB����v�1��Ph&��r~��:�_ɭ����k��a�r|I��+gu����E������#�A�7�,oE�9c�Y83.2�I�)���D�@�3�1UדEG�J(�ex�&���G��S��.Q�0� �س;�?qD���Y�8����~W8f>����Z�pvk3�|�(���OX�b����q���M�6�F��{�*p?c��V�Z枍���2����8����������b��Ϗ��|8�l�Q)>�J���;bL?Q�H�S]���Ć��qՏ8�j��]���k�|T[��a�9d�o�"s��uJ���3(���E�Z�
�%	�#�.��MK��&���5�|�*�@�2�ޥ}KL��<��**?�M, pӄ�Fc����!�k���<)�_*НfCj��>��v0�4q��b�'5Ԭ!��S�~���
ǟ7���zf<q��辦j>>�KѼf��'�ΩS7r��qE�]��N�T��} z��ـ}6TR��.�г ��5g�·<�Ľj�sȠZ��̶Q�~�X����mk�7 �g3%h.��$Mks�~ܓ��<�^ʹ��-Z��nf �r��k�տx^�λ�j��I��Y�v��֏Հ9�	s�]r�8n��[�._��5\���A{�gI'I����
+�4dC&��w@��QuMɓ��קN�����چ���o�#�yO���7���o�L��`Y�)@�j�	��: z�EM�xiwc _(��`��L�>��wq��5r��ր%Ѫo�Ӱ��[�Z۠��W�E�к�W�_��ws�F����ۈw�`���r�:�6�ׅr�Epd�pR�:�sQx�Y����|���@��Ӱ��q��R<�#�q�K:�t����6���ɺs��3�$�p��\؇Mr;�����Z�w��۬DC��A\�`��H���uQ�SB�@�]�+&�O�/	������ړ܄5K��<[�ZC��`o��'����p�5UĠI���A��p�KT+����߉%"RC�mzkZ�#�E5#]'	$K�3q�s�T�m����q����F���+H"�t���;�L	�C h6`�XI�������f�>]՝'�>d����G�M�y�!i'29��/��g�W3Xl�?�`#
�Qh���Er��׻�A�}�~=)}�Sj{�,���|���#Pk��,+U��`m�e�m�:/6��ֵ�h8�	�٣W?�.Ñ�E+�i8V:�L�ٳԬ�1���N��J�.�heA㡐63Ǫ��)0�P�4�D�%%DLTV.��q�̅�z�:]d��i��y�	�0��M��bt�b��B1㾶 g�OW5Q�r5W�+י7�'lN]��<��N�k-ԙ�^�@�ԅ��S@?�z3�S�8���<wdg�S7P���Y_H�b�����,z$�_���쏵*�����������E���h�8ެ����8{���e��m�"Z�im�P����PN��Jrw�1`�����_�K(/�r����8��˱�����H�$9�W<�������D�bTYD�"ʉ<�!�H�������`��mC���0�a�"sV�a ]�G�o�:#;���,*;��]W�w��B�y����>�W��W��\	b(�) � �DY��<�`#��ɴ�n%v��x&�9(��@��T�i¤���=����(��{iK�~�t�B.R������1x Or�Ȓ�*6ƁU��/+
�@��is�&\�z��)XI<
���W�B0�@��%��hʌ�Z�+�G?oC,*g�����u��}`ʦw���{+��R�Nm�:YbZ$���**9Nyd#�U���������3W�2m|�Ƥ]��ں�8\���0zɧ�� CI�q��|�&�xaV�����l�W��@2�����އJ�hƼtFO����F/?�K��>}�I���f�o_ڣ�LY�h%Y�dE�tAJ�������ve�DI1�0_��#����]	][hH2�x�����iQ��QlrK�X�}H�jQK�:�Y�*q#��tu�YB���c�dZ4���A�@Cc�jqLz@�E�"
$�v<GW����U�*1p�ᧉլT˞pO�ڃN�,
 L����&K����\�8�P��v��[rL1mSe�,�*c�֤��R�7!䝵8�^[Bz�+�u��U<���'�8���9A�I���s#5����(q�=ss>Z�Z@~u�{J��/+U�kE]���d���Y������1-��*XH���:�63#�̿����6��>��(� � �lN�^��h&"��ޑ}ONR ��<'͟��z=���$P���ȕ я�Ԟ�.�u�q����5D��ƣ��\�*āّ�×&�O�K��u�&��k�}�|�v�;��=� U���=n�[b�b�N��ږ���=�ic��v*~b��������Y��O��ۤM�
�k���*�V�Ӏ���=�6�O�`�Y�r
 ��A��՛7�c��{>�ƚ�L��c�Y�J�&A>jcx�͵ȑ���v���8���H���Ee���>��>Dfh�
�<[�oR��EĲ^�eC�?��Zr��uѸ6eNK7�q%�5`�d�i�`�%V�}oP���g�;��$3�+�i�@lPy�7FN�5v��W��ժ0-K�}7�K� w�i��R��O�;�J.EB8e��O<�W���}���Zk, [Gu�����1eY��\�W,���HW����}�?���
l����xf,r���:4�v?��S�/�
�ЃE�&A��OMI���$-�����zI�O5RA�I�uk�ײ�l�\����BHO��g2����f2�H�������r3�|L6��$.��"��s?�4��Jƫ(�rI�>�<����~�� ���$S��(�+�"�y���������pb�aO�t֩Cs/v������ב��V��S�/.o`��ޙ��|{9]1*��J�:Hh�V��^�N'�a���+��"k�������5Y%~,�J�G�uVc�u���m�25�IM�B&a�f���Gi�8��UPd�<R����:�"�a����I"A����s�����*�G����ў�=�0��'c��NM�|��ߚ���O���A��'�SԦrw�r��������n�(�#<�\"�������)/�W��WT��/�olsF�~.�W/�A���S鬆L	�A�m��	2vV&��$p`�G�:��N3P�����������G�*ܪ�٣i	���k�p��C�����D {�-ϐ���E>��Q+���Q��_g��ȦT䌽��a�s.p��l*�����v����U�X��kFZĩVin���ڑ�c�EDV�t��82>ÀA1��R�&�i�iT�z��*i�)��$��H(�*�����zU���Khd�|U����l_�߈���4�a,�N�%�8v'  ���
�v��(�:�\-j��3�� �b�}xp�1��Q�~����_���=��{��hMaUc�P][�1� tgƃm+[zA~�D�ɛ.��u�Ԭ�:Mw�)���I4�3�D0���o�ZT�*��|�,wU�l�a�t�@�.�[#z(a/d��1E�z���z��GgU����̗�k���&��T�:N~4!Z��D|�獵t�W�-j�R�GǕ<�B�Zo�l\�$��q.�s;!ݠuu��J��w?]3[����7��U�:�����;�*�T�U(d4�"[�Z���j��gE�'N�!|��d��������p�D~@<��+*۝.,�ػ���Q(�Ⱦ9��=FF:�˟j�|]tT�$1cU�p	a?�.�###�kn��9�-��F]:):�����#��λ��liC�ڴtL�;Xh)j=����B�zߜ�E��gh�m�'#�ҧ')�};E�r���Kp���%��S�nY�ȅWE7�~���%\�avڌ�y�\�U�]�C�{`o�g~����H�n־i"]y�y�V�R�=�p�h��E�m|��x��y���wl��_�/����D�W�J�]^�ʲ�2�����&�zm&�[S�oT�f�#��S0oٹ�WW���^C��5tA���1H�n7M���Zk$���^_�0��Y+9��q������:̅�92Y?9�j`���X�M-/@�b��T7=��	ƨf��m�t�.k%��9o�O�)��0s����!s��9v������׀ ����{�����X�ŭѱ؃x �1�ۏ5|P�xݎ�Ux;�m1v���4��kp�L*?q-����\ʆ 6��2�Y.��SKcu2z���F#Yk�}�t�qB[&ݟ��h�Q0d宦=�F����~A�2Rh%$���3\��;�*Ti�b�A��%�0�����3I�>5��
���JՂ��H]��W�U��J!��H���g�;��@|���9����?B�W��y���(i�zZSFBz�ϡ����_=IwTj���=V�����P���&>.2��y���޺���H�=��xz㩯��(�O���`:��2��B�-�1X5Gw.f�;��S�G8���ÑW�]L���a�	��(P�-�e�C^���Ϲ�!r�|������<�LvPoN��Nu�����h���`V�K��Т���p�v���B�Vc��٦ATbŢl%�Ҧ���V�c�5��Ԡ#��t{��4e����L�>���`t$��P�:�GI<=����X"��1�@�,����5X�3Q<���+�B�j�����3+˸�%
��2�U�ps����K��V���B����Gs�ՠU���J���+KW286�����8%rj�T7����d�����Y�FR�����'d��f��e=�7&O�Slխ�!5�%�¦��Of�}��=�<2����B4�?t-����*��&/���l+����;�����vb�`�	���Fm����X٘s�N2�|�!]���H��-�����'[���Y��Nq�B�z��U$��C�}]ӭ���=�Y��6�U���мb���;}"�#�6zJ��c��ʬΛ�x;��O��д��_(B��4�Bg��qmmd�ɪ/�>NDA�|.R�D��g����_&�X��C�l���I�����5G�~f�PF�}�W��զ"d�31��p4��g{��zA�sM8�8RKA�+���LS��P�e����oޯ����E<O�@�J����:~��cH�����&c}v΁�M�*Y�Y
ږe�o�=�߼��v,��魴T�\(��y�
ւ=m��C���h�����B��k��PVK���@�ͼB�F︋unX�6�@G�/ ��mP=eM.uI+��w?�[})�cN�'��������6��8��QDS�z
��ǈ�D��1�M��s4�ge0z�:Կ���E'R��<+�`�{��ˏo���L�擙\솢D�@L ���Xzg?N�`ٺaԕ��@Ņ[f珚�;.�s �C�_��UD�[���1|�
gd_���!�j�s����!D�s{K�u��A��" �8�,P�_&�(�D�&����e��_���d���?5;�D����~`�]�Q��87�ݮ&K ���o=��Yk�����V�J���\"~&��H�N|28;�@�4�
p�o���oD���L�m\���k7p٘$ZB �b����$����]�#��ٻ�W��x#s����ʩ�̄g���0bb�BM���5,���7�6U��V��x��
z��~�vq`�p�H��D?��2����}yM�e�e#�+�:�2�35(ȫ����m�u�ֶ'�`�t�����Tp'�?�֏r�h��r�-�2S��ߑ]9t�?Z�dK�L�Q�
+�ϣ~q�!��)V����b}!�t�07�ğv/�$�}����ذ(��zXn���:���=��mX`�n���F��@�F;���m�5{|Q]D�+���� 2����h֔��(3|��l�����)_ ��֖Ku���7�h�)�i����S�m�7�9P�q2��r�ѷ$�8�$"i$N��Q�.�@��G�˵(���q)بMh&{�u)��7.��B6��	�q��l9����؁��&���;0d/ U� 5�f�o��!>Rc6z/�C=i�a�6 ��~do�ˎF�+��"fD�?��5ڑ�'�s�����������c7*�z��7�=.p>D����J����״-/�)6t�{�{�>��aK3u �LZ�V��Ҧqi��;� \������xk;-����|�,�����yC�:$Pݢ�0R&���Ę��'�+�� �%��x8��G�3���mBY�1�������{�(A�������q�ˊU�bb�b(7�$I�V����j��5˂*W�PX.7�,�d�FJ�0�گc=+��5
��C4�Qr�O��Wc��#�#�Q<���H�F�@B�j���В~5��X|��-�;�'�e�CU+�TP`8�A�c�t���
�jH�u͚�,y�Ӗ���i���r|)���I�9�L�"w��"�[jK��{�j_�S��r��b����e�n���5k�"~���0f����� 4Xc�Y��:��,��pJ�y3P�@����?.z�vF�G�1��6ʎ��D��ù�֎p�9��oo\}rJ����&�T�1|C�o�lчge?�l�4B���ד^�#>���n�G������:5Y���|�xo
l`r��V��vpe�$�uV�t�"�C1P���Ǥ���53Xm�?*cuY�X�K�I��� :���g��@qu~��鷧)�:�\Yyo�d�F�EŐ�Ek���P%<��u���&��x2�~.��~�M�7(�=<��)$aт@��R��W���(��.��C�Ց��;A�X��1xT�Ff��a�Q��9r'#yi9�:�l���� UG �d�\�IP�"�� Z�~(������ED9�̬e��@1��H�a�vd��t+^�O��G[��@P��}I[Gf4u�ja����x�V���҆[ډ�QFv�T��*����{ɥ��Y�>Ł�j�s�Me�o�Π��͂Z${=a�qW�-h�:��5CC<�+�\��nq�\kKar۶�Z �yr�0P���)�Ib����VJ�P�+�S,_�c�N	�:���U��9z������i��\�m�/�J���eO���H�[^yb�v�퓰RΊ�c)��ց�S���8mT(�?�~@Jݿ5Ϥ�����|�[S�����	sv���3]M���KX��,O1�To������<��VE�o:N�a���&VH	qT0�`��f����R56��TSʷ�D�p��+�A��d��4�AV/O �����V�`)adm��Ɔ�3�>UH..݃Ӻ�Be|�0�ZF)�x�c�_e����wԧO�?N���0CT��|��j�(!��qaX�k���?x`(�CYOl���-���q����ŤcU4�q���gMދ��7�G�ə��a���i�V�3�+��"���Za-v����_+���Ҷ���3����MH����YA\�`���i�'�_B+����q���y?��}d'/ʃ6�5�줁�j����ҍp�ص��,��W� =��\�E���O	("|�ڟ;Wa�?ꙕ5x!`���W�w��&$F��V��-�,Xy��] �2N�B(�T���z�xR�$e�3�(m�+��ơ���7ԉ��Q�=r��V~�u3�/�^���+4$`��dM<s����Vׂa��>!K*$aP^�$l%K��A���y�#��>�}-��)h���բ�EE^�	�E�����F�oAX���$�����BQ������+K�`����D��������ݦ��a��b���[�(/��%g�%�xH�i���KY��R�ft��Wo����3�?PBnΣ[>on��^PP	9�q�#�s�Dy~�Y���6�m�S���Idf'a+�^���Y���z�R_�BN������`����N�
��j�[o������1�d��3^�81���9pd��Es�����QdĆ��H]\Sb�T����f�Z�?�c�_46΂h5��E�X�����Pҳ��̔$k����,�(mOi/�k���c3�>�my����	`�7{�z�d�ߎ����nC�����A?�����ڍ�~�(Ir�d�1�'HJ�>���)�sƵN	j{� W=��SI��ݿģ���74j�xTh4���}�x[z,NF�1�}��z ��xȭȭ�`iP��f�f|�a^n�����X����ܽ "�����m_뀬V����6B��#��i���%��	��劲;W5i��oO�%�A��{ɺ_ �u�d��T{��i�kԥYy�ݰ.����K�}	�ժ�;pw&�4�H��<@�PD���DxMÐ��k�jSۺ$@�
7����s;�;�C$�m`_Y��T�B�G�;��ؤ��e��kKp^꜎&T���V���Hh�n����7u�{���:�][��bS��L�5�{p�s��Ɖ�Ԉ:ހ�H��3�E�1N(-�}5�R��:��n��n�y�k�i��d#ؐ�CC�K�a�H���
��I~2"�n�_=I��S:��c筞ui��q�?ğ� ��R�^�k�D���Fi�T1]�+x/0�U��jB.�]�~5�eӬ����>���|T\�2��~n�~���$x�0�e����EP�N���,4���Dܹ�
$�d\	�*�U��뎍����#z|�{Q�c�E����V���y�خ������&+5�&��i��|C�/�m���".��Z��>D2�#�R_�Ig_��pO�ʮ���2��}fM濶��̓����?a�Uh.0"��b�Ch!yY-�@ �rS�G̘�s�˕�9�H��uœm�tEy�%��k�/M� OG�ѽ�l Q�3a
���\�b��0㲈waTk]�5��.6��N��������x�V�.�P	�ٕ�1�v1z��9�νxVlc�E���D��Ve����e���<�Pwmн�
o�P��u'n�	�E�sG���ј�U���.�yf��Xz��u<��I�P��<ϲ��dH�`
��?�4�)�jsXw�ux\�{:�g��IŖ���7+�X��ߢ�UU΁ER[j���O��[E���,Ǉ$/�Z�gp�	��A����9����<,��:���1E���+|l�Ȗ7�iܳ��iC/m&n�"P*9�Oʹ�Ct��l��g\�d�N�%���<�6/�u-[�E@X���ݽ�S��с� %���9L�%Rԙf�'8�>,a�ӳ��<W�?��|�L�ͤ��8�:L���>��W��L/-e�a#t����vI��U��R���+7hS����l�����h� �^� Ԕ#���d���i�&��Ú��ӹ�+�ry]`s�Q_/�E	S#	�m��\�FU����)cW����u����
+��G3��:ūwT�4���=v�(+�ʛa]�ϡ�!E�-A�WL��M�9_Q����	��8ؠ5}��;��,�����*�%�b��#1n��'i/�<�˷7��H�������Q���B(��+w��C��s�&:��XT0xAntƨ�;�::���X��������E�<]<g�q��Mn��K>�<����7�ч�����������n��}F��o�NC��ɓx�)��˲�xM.w[?W�%ה����p�d!�(���*R>��u��C��G��o���<uY���m���5�O$��!'�&�2Og�&3���~RqZ�:bAp�����B�������1 �2�®{^�u{%���*ۘh�	����E�=�@7>o�oX��7���a8�.P�w��a��@����@�=F�1.L~�3(>�!��wl�]U���p�'���5����ᛎ�V��*��}�u(���v��n�F��t̀/�O'm#b".@.��Rv֣ʉ|�@�rjƹkp�wg	��:C�0���bp�à��X�h�
�b���n�=�װ�q��W~��E�|I�%��ծe@����X�?(P�0�í6~&�����b�w3����!@�f�G/	OC]� ^d�ñ_���rK�(��W'=�1�зȐ%������T�/=������F{CPԓ	����9�K��hT�8�TM�"y���Zؤ�-e���k?gɮ�Qȝ,���!U��`�`o�K��W���@��4k�/�'�V�^����U�hQg�� �3Մ���.�Ds��Jt���?�<K�vN���5�F-����@X���u��&P�̖�,��"A�c���֚���q|	����q�u�q��Oc��)8�S�5s4����6��N�М���Ӫ���-Q���0{A, �^c����'�X�LD}�K���٬���>)	fl�����
�a�#�2���V�+b�Iol��zkL���/h�P��BK&��a��[���/���69rM��{�aݹ�߱BU���g-�	T+��:���$�ϸ�ٯb�Na�����^���Y��W�x��(↪��4r�f�/�]p�:�W6��#�*3����t/��b}.�<:�Ԝ>��i��;�Θ؄�c��荙5�уI��)tO��g����l�K�Wj>��%����vIE�f�t����1��=�-�c��㭬��vkԞvdGw�)����0pq-�=o��rX:�<�#���XW��XLՋv;�<>F���$֎V�Ah딚�%��[LP�m�5W��r�kBr=�6��6����lut�ˠޢ+�$Ppzkv�97N0���!â�$8[����;��1O���VJ�f������Tl��ȇetƲ*T�h�`��R,�}"F�b#*N���W�~@ힻ���q���W�k>7���O>���,�2�wLQ:xw5W^?/N�m��^��ރ�]�%�:���3g��t�e7�O����c�6�(p$Hn�3]A�|�t�ǳ*�E��,�ޭ������ś�Ȳ���.�v�ṦS�;bg��~t�ֿ_��7SE�����2�9?1��%��n沲p���PU"��+Hj�B^� �
��AR�)l��K��MD�����\�P:o^7'KdGv����b� ���a�2��>K����p�9_�w5�����kyLS�A;W�J��g,�9�gӯ�:5��2�|��$�.h��>����зnj�.�7צe�2z�?��0c�D��D��G��%�=Σ(�g�0����B(�.O�׀y����G���c=��F�+��6���l��Fߴ�-{昖��c��6�0xڏ>#����"��;r���J�'T���i������+��ϼ�
U��~��N�����D]4;m�~��Nՙ�hb�)�F~���l� �h�Ʃ�;�x(�ѣ�<������bt��3�D�^��[08P��Ԟ`My��j�~���SP��1�wA{��|���cM��׶<tE��nQQ�.D�]�>�\�']>?۔�!���k��;�}{�l�æ�RX�\���$�5nX�����Z�[�g%v����Yl%^� oѕ'f�R`&�Kd�~���E����Vzivo��jp�/��%�+p_�ATN?n�o�<;]{���
V\�$=�-_.W�F8�,�H�d���iwttr�d��gx��/�!�5y��Vj5��A��Lw�{��T����?�1.�T�fv����*"�e�ł���=���jy���O!%}�6�t�{Ou@SE�&�ØZ#����ed �x5���⹓�4ڀ��t�`���Vv��#nl	�~��dӅ;���������0�M�q�%�@]�f6׊�U�B�l����]���28�ů`}dL�A�Ϗu�9W����)\���a+
͛+U7)��!����f%�4���H�ϭ�)K�����U��Y1Į���\n:0��4���l�l爘�y�BY���~H�V﹬e�V� ��	��S�_�b���=��[E2��L�ʫ6b$����dH@�zV��UA���<����2���j#蔯?p��\�2�Ui���þ�n�����PG� (L�h��fq�m�NUR��+R0W`9��<,�{������J<+�LI(�J�uzV6ϧ ���*:	�8���oPf&g��)���0����k:�?NT����wE7�{7yC�:��+�[s�	ƤOm�c�ja�����;�w]7�ч7V �܁�����5
m�-mBN��-u�_��m%�|�(>u����F{��O�SMpp��M�o��e�ٺ-	8l��uY`�4��{��|7�H�:#��;���D�*���4�k�W��&����pQ4�ʡa�7'�3�1��{ʏ�C��HFX�v���b덽�HB��BO<�
��3\�C��ɣ�}+�t�G���.���A�4�*��^�܋��P��W���52��'H�5X�R�v�?n����]�,H����q|������G	/�
W�K��$�b5���$�=6U&�v�0�D��d�H8��*ۥ~�W��f� B���� �Rz��KԮ�Do��ˤ�jm�l͞�,L�����t��;�f-ᰆ�ڤ���7�L��A�	cӲ(ʰ(�0�n"K1�2 X��u�KdU뿪�8�Ԝ���oX�����./	��g�����������o.Y2x)���#�`E&̸P!�<d��!w+�����H�u�B�N�3J;�=oQ%�Qq�WAYB��h�؜��N�ڀr���E^� U�҅2&���e��)]�C�����:�䓉�q��DI�1�V����78��V��/8
�S�f�d ���o'�3:R�$
�W�m"[���~& �Clht S���q��I˅H�|4���
%ȝ�i.Kg.�_�p�|z�Q��M�Z�Jo�'�� �8*���V(t8�s'tS��xx��������.�i�����.���Y�!ײiޖm|7�S��p��Ӊ2#,q\����> �]�\���%�J$7��ŕ�{���+�2������=J��[����ј�� �ƫV���c,�t�?����I$ �U)�:�K�^�S���,iA�7}򎟸4p72/�b��t��!�6h���*���s�J�sk�!qh����vS�tc6�R�B����x�#��yiH�����o� O~z���9�:�e6ߕꉃODs�n�����Sۄ5���&����v��h��������ή^1���`$�U�ONX�c��+Q�D�X�ڱ��b�%�������В���v����t���̴{��\h���D����H��J��
��@�}qk5N{XT�kK�Gk�ŘK컸����简a�+µ����x�n�k�FkJ��d�6b��p�ރc��κ��!����	|1a����R.�.�h���'���:�Y���|�>jҢ �e�?�4ܑ�`2��{�T��w�`��D��g�;���X*�.�9��4	��iV��Cn�c�aCyZ�<��Y.P�zD�<�gE�+����_=��I��v�{͔4P�R軅������T��� ��4>�uN�ߘw��X��/�j�oP!=�*���^f8�a"X�q�%@�}�@+<��2���S��(�]�y�Fn���&p��V��R6�;�'۵Z�ގ�hUΝ���~cs��������hK�,rlz��1g�/����\��ٴp��`�0MN�'<��AbS?9�׉���xs�g;��T���$b�pL#_c�	||D���ܶ�ь�(�c��\���2G<���%���ƦM�'�%L?�� 争8?a�������B��b���\z�(� a'^� \�_A�5����g7�!��>�2���˝?�=�J̏����'�<@^����f��ʞ���O��x1�C�G��]���ߘx���ST�j��Y��$!i6&h�Z�O� v,n����Ss�U��wf���j����d��&&]������<=�B�ћs�NF�e�l=�w����H�_��ɴ����p��F�Lll�YP�a{rNID�=�7��Q
�
�5�=;N�~ʥh�,��e�)������bI@����Y5�n��o�D&)�b�<���⹓��^IwJJ~z��/Bh�{#��� �`x��V��k%�A������o˝��]8{�t��# �W(	HY�쥅;��1�����;�pޓ�M�&��M�o��s��=,a��v/�P�:3z��������M��eԘM��w������N9O����|�!�CEXw�tw���Yi��;�8��s\����lE]���l��x�Mg����L��@��4�:��[��E� d	�����!_����҈�[`��BH�Ym��~���֢$��_I�����`m��2��TÕ�����ْi�^gYiK�ԿY�x���	�y�T:�L]��S	Y��k5����3t��=|'��95ɝe��x��mb�`�_���%��c�F+��J�mJ0s�xk��%4/#S+ڙɇ��cjpʹ�7H@&�dv?�����cj�"e����tU�9g�!���6tI�.�	;���)qۓZ,��8+c�8���O&�.�A���N;{�p����*V�_3�l���{��t��R�֝��%��V0we�p���:��Q�����1�%ȷ�x�
���u�1��Ҕ7	g.���Yv���Cs��ћ����j+��T��r�-��>�����@��	[�Ckcۅ�&�b�ci�#l&A�l�]��r��)J����S#2ù��w����_�洼�O�˛D���#nr�(�E4T!K�03�����m*��h�C���d�3�7g'a�~��.��w8,֪�8Z��ã�x
�&{���wU������^��M�Q�ů��g���	��j\R�K�(0_j+r	(75X��K&�r�� \Ist0�Lp�3�3��o1f|S/'��,�(Zw%���E����$�j9]Fx\���UY#�����y�ޠ[�h9�qS@�����!�����c�]�l�%2�/R�7� ���$7dR5�W]��m���ŉ��0,a���V3#!+4��=��/)?)#���2����	�4hv�f�X�u�YMx�md��:Y	�`��h���6<�~�i�˒;��Ƞs�՛90��
�[Ŝ��֏��������_[g�ÿ�q�\���5�E2�P|�sS!�$���7��a��=�'�ʻ�ۧ����<��۰-7��<��z*��,H�}K����W�ݨ�y��t&�NA)����K:���@�oT�W�����!oٗ��gy��L�®��6rd�1����Y�F�\��W�䳟�L��U���C��a�"��k�Ɵj?�?���K}O\��_h��D0n��.\�P�x��q,���Y�۷i���ٲv���������J����d�kpOԆ�.�<V�p���o�q�%n5jo ���Y���f���(��c�ct��0�ja_���#��U�Ȉ(-��ڣ6-��r�c��W�2T֩E��\����[%���i��e��v$��J��e�p��k�4�Z�34J�:ѹĴf��Ҟ�i0��+��f�S�R}[��N���2>L��I��f���^�ޫg���q��$�CFl�ߓ��O?LT��Y.���s�zIr��LE9y�����>hހ�2^�=j�A1�g)��2���{�ڜҲ�|���'Ο�j	`�qRn��ͩ(]�p�G�XW�+��e��	�Q��o����0}g�<��j�E�Y:i�7J[a�Sc`AEA�����@rozmH�>�اe}Gb��	i0�3k�r�D�vr��|3̠�l�Hq�<������aM�Iiѭ�v�Z��mw#ևW[���=�\\"5I	��� ��J�tڊ�W� h2��;�.!d�ǜ�M�=����Л�G�|裸�d�0�D�U�=�U�eH�o�Qdb6���J%'��ax�(f�$V��oY��M���z�8@i5�`:�z&����[�Bԑ*����=����;�ι�u��=#z=N��s5Ct�B�;�4��G��1��SbӤb��-�P�O|.�b�VN����|���*���b��w��(Kz�(!Y7"��a��1������;�&N�J&E���J8��TqfO�� ��I��]xT<V���c*M��t��O�#��q^��������蔐���9��e��E��5fN��!k�Y"�ōDQ���*m�e�[ �Ί]Dfj�1�>@��-������&y��[XBsh��k��k0V���1�~X+A�����EL�q����a����dT���?'��cX-�����o��M&(Ձ8�2a4j�4X�z�?��AJ��c�޺N�����Gs��>��yo�iUNܽ���hL3��k��ۋ�Ӏ&�⡔a���ٯ2������5�
��<�6�(���0�ƚd#�W+�~����s��t��(#؈�>�fq�|�%>ڃu�f)��� 7|�	�?i	}+� ���0mx��7mŘ+�%pb��חb��p��w�9�۩�u��{k���K�����a�m����`O�+�8�$�iP^|�a:�\����R����0��U|�U���s�y&��o�{��}n[��<'�gw��l����.ۿ��#>�6�W[���N˥����(��>�^9(�Y��T�J�熘��8 �z!I�t���\*��s���,��@_J`����q�۳Fq��˭G�^�!qR_a9�%l�AN@�J�@��(��o��>�Gtj��p��p��X�s�V��fU>=>��%���]�Ci�S dG�Q(��x,�N���Ǧ2�`��o�S����r��[D'�4���dH�*t <<�h+�N�ۏMo$��d�Νdd�#j��j������R;�ż�y����A2��rt�'Sg�Ky༆��'���=N3P�U��D�1p�Q�_�m�pŬ��;PvtS��� ����j���'��#ϒ�~گ����������%��}�l�?�tf�j�,z<ّWQp�i[�]����b^e5'A����ⶈ���M�=��KVQ��X>6�����E��bt�8ڟ?��f�h{�"<5@ª�pr��:����D!��.+!V��d���01��n�̳��P1/������X���~�о�w��\WW���g�����h��k��}�.$�eM�yr�������}�r�CR�Y_�S�7�HI�` b�|@w-X��|e� ���>����I�5��kMSU �</�0���I�m�\!��U �&@F��_�ba�9ΰ�├�(�1<:����(Q�΁��s��J$�jM%���^s�%���)%	�DH�PE`N�lea����d&�R�3?;�����#���Փn���|���.���� 8ޤ9���M��!p� �ƈ�d�ga��؛�Q����i��][���E�V�ز�>bt^�%t|�͔`m�W���PR�$���zr�,�J$}헬�*�u��mj-�s*�ɀ��-G�C����ଃU&1=��E����F���3�� �?$y���5�A`�vS;�L�n�`X�6�7���s?7Ǖ�n]���B�އ�J�UQr����߉���Ligy�f�OOB�1[Ҝ����cUI�J���5<._s�P��ٰ[������/��4�C�ct<Tr�Zūo0��#��U"dU�̴�`�]��1h������:Q�Fe�"�u�7�9U"#@^��o�Yk,��K �{�s��|���S���j�=a_.�����M���[��g����'1ϐ{%6B)ޅ<)S��]��Ƅ��bn�*�v@������m�i�D��@�l���3fyv��� ��-�p��8�n]�z�/�E	�w!:�վMp�r�=w��t8��!��}��s�v�Ό��랰��Ϩ#����B�����B|܎÷��ԑ໫�!�GVFc),��E�ψޜ꨹��V%AZ��K�$̜n�o`��2�u�50�`���rӯ��#��M�V>��f-��LW=su�A��l�#�.)s��~V�]!c�S�!�,�'�:�}�p ���fe�A�Õ2owZ^��X%��UEH�N�����k'2!t���~4��x |��f����=$��� �^U�-M�̳���&��.Na�w&?���0��{��Qj\s�$A���揂%o�cfz`�m��+�e�3F㮱S���[�$ �n9a��Ș}���(���hWKi,b(�i<�
G+fC��K���8���@���
Ӷ�)��#m>a���g�$(Fo��p��.�<d��ѱiT����wb ������L��^��ec?]�My�XJ��c����y�z��u��wɄ}��bEm}g���+�ξ`�þ�
�mwu�z.6?J&Go���p�#,@��e>��$��e���y=Z1Ynd��/�jd������w]�i�xC�c|=���K��W�s��bii��5�!�+*�q�UF��� �T>(Wq�H����t�ܞ�6[�$��?�(�^�4YT����Ɂ�hL=�G4�� �tZ���M�U�$�|� ��Ȍ���J@΍�p+��O�W�fZ��;��B��\�D��,*�To��F�CŐ�Z�<1���7��硤N�"����D8���fa��e�ȴ	O�����o?����K�X/�ݑ��ßb,r:�����h����7�O��2�����<8���-���8I@����1w>�ʆ�:�5N>4�L��z���ش�f\��T�.|�������ίn7Dh<�����$t�=�,�]C9k�|�{��t�Π�в�*�;Q:Ae�d�� I0E��m�˧A��y=ɣ�~BͨH6�x��0�����ҋ��  |z_�&�f�0�,4Q����Y� Em-�8�9��[x��@2�f�w#A�����G����� b�4F��3�k8�R������"�V��J>�L$�|bS�gm�y�0h��uM���&h�=i链�,��E����'�Ya���g��\ �O� ���졁�Qį�ly�8�n=7��i��������A��F]A �l��:1�l�9=n���0�h/G}̈w�D�'K��9+_5�Q�=��J�1	*@`���$���1ٍt�$�\�̈́�e�׼ݬ[Bf�����[��^-1���N��"h��4���S"����К�� j# M�ɩ�##.-�7�+;T%B�iD��v�Xd�����Z��M~��+E�m_�h4@_D��-z��&8�N�	.ֵ��J v�vHݨ�`�ݙ?�����g�����S0�I�2��;/w�-�Űэ�9������p~�k��g֛�2�vSN4�}�y��v^����Z�N���<C���S�,��J���g�pP+"�=끏��"�T$�����u�Mo���:R搭i�]����T��/�{%Eަ��p-͑��Uϐ�8&Y��n"�R�p�I7�6vY�'U�@�m�8d�#���� P�+��y�b�X��b}R���7K� s�e^��9�'yC5y�:�����ixO��n��x�}��͉�_P��������~B0\�[�J# �q�l�<��z~�Fq�DƇ@�	��0ce�9�$���v����P�Ά��P�K��O+�/���W(�����N�2�怒Ȩ�I�?/���-U:j�;=E A��L�,^I���)�G���8�>Be�}u��Oy��'�4=rf9�ט��/Ѩ*@ �A�BT�%�;�\�� ��N�Ո~���GC'R��	Ę	��rk/���'O4i���~����@�`����5B��0]V����J�6m؄i�
�f�	�#��Eߡ�b����kȃ���d�|H���xm��5%��LHQ�� ���drFFώH��j��m�:1�+ޗ��W�4�DV��j�&H���EA����5�S�`�{�C�s��||��j��'��c^�@��֦gڴu��G|����g��X(U;uN:�_��� �E���yzi�C�?1� �D�S]{��Y�b0=n�B-�g���<�܃x>�����z6��"&��t¼�Ne�Wq^7�Y?Ӥ���-2�re�	K�Zi؞�2 ���r����L�W��d����y|�a�I2|/d2�g×�^����p�"&/�m�"��ؖ������)D�c���ۏ~{6�'��:�����h�o�_.L@칡��Q(H.#~���<���!��Wo�>���2��@~�'������ke��g���[�%_my%l+��e74n˩�	g'�uz�R��!n|�:-Qܤ�^	�
�Q�͌�z�c�P��eE�#�G�(��ٰ��N��W.���↰V�LwM�X�_3IH��]�/ �`�z
{Y	��<F���Eꉕ����O��Ns��6��|�5���Ј��6R<��M;�?Z��h���- i�o|Ʀm�;�א�M��k�6�S�0���H���?y[t9�-�~���0|F���g�i\O�UD����;�r%��xv^�"�I���ݗ���K����_��bŒ�ei��By��8"A� :��,�M���@�[�b�]O8�y��������	Sn��.�p3���-�����B���4Wn���>��3e�*r�+�����#%��9��`��h�}z�T����pxD-<.@�J��́���E3�J�(X�'��$����:��a..�uU�띄$rtl5�
�_�C����2�Ҁ3���9W�'ke}�]�[`n�pv�.ĐJ.������<i'SEC�w�H��N�����E�_E�.���~1��09�p����BUgC`�R�'�f��-��'U6X<e���B���)"xXD[��܇���=iV*͛1�[�|������8�Z�"`N��'i
�ta� h�W���B�?��oAj���t,���W�n-l���3���-^���O�ݬ�_H"��#��j�:9��`�hǄg����F�wB�DH����W���d9C_��Ke-�o�<��&	Ix��A�k[ ��7�Q��C����&I���^9.���,h�K?��� ���$�%�D���[�o�Ni��ypY�	�籟�|�X�p����$G�xK�;ۆ:	:��Q�|�/�y����:�b|�#������~_Ɛ0��+`f`D#c���a�$5���µ{s�s��D$w�ne�CkhUe�*�wj���n�8�Er���5�*]<�P�#�pk�X����h-�A�+���:/(��!��_�j���7e㔽��haU��#��=E��� GQh*���j�,'��GG�	|t�U�5�Ot��@O�!L�@��pA���{��sE�ڑ��:2��q�Knbs>@�l�̴��0<�3��p���B�����������o2i�~3G���n�bVg���.��#�h1��l�7��s
���9OTT6�?e��v��\�<�B��;2� �o��.�xWvkWFu��C��������y�Qh� ���co �{�xQՕ�g��EJ%��.�XԔe�t�a �y	1�^�D��riΥ��T�����T*Hz����V�Y�w�(ˎ�k����Nq���齗}]�U�#�X,ϔ)b�t>�Ce���7t�c�*��i��J��l5o�
x�I�-�����q<� ֙�G(�Y������D& �w*�Rt�n��vl��n���+VAu�I�E�!�����e�ߺР%>�\XԖ�h���oiB"r��������ܶW?�G�C'��ȹ��"VcpYVB��m2��	2���%�ӳ�q5�_W��Ak�h�!4O7���n~߮]��o��u��ۭ��-�"���[��^���A�6Zt}��cP"�Ɲ ���W�Ncy���4�.9K�+�����B��E�;t�{(jWS�0��eE1T�X���0���p�W��O�;X@� �P�T5&�:��t��X����~h�%sU,�e~�����}�h͛p%�ꩍ�$ʫ�?�F ��ڍw���σ�%�z2c�:��5�����E2 �d�g� uQ� �*�p�%��Zp�u�?J���X�T^�� �-ݱA�Wl,�Ze��X�C���T��c_}��;�0�i�Q`���q>�r����ă�5B66`7���N��m�ã �t
2˒[�П{�H��.�IP�S>'}u���]RT۷ ͽ5��CVBWnj�&���a_���ejXBzt�5�{�ZIBY!hK#a�x�/��q�n�8ɈZv�i~2�'*u���A�_�qCb7b}ph
mĭPgq�op��^�T_��ϨI�� U�'�x�S}UB�:��*0L�1�uu����e�׾�A��Xg��\��@�ޖ53��Y*����w���f0�1о�J\ϙM��[���^�����;�򗤤y;��
$�xP�#�W���P��i5I���;!�WQ� TF�ZI�LC�{^Mq�a�%�i�����x]1�Ʊ?���\�i8DVd�'_y����Md���z����^2g��`p�Y]a[��e5�Op��.ed�%4�B�?�*"rs��g�B�;�͓/j?�	�;=�N�H��y7�Q�'���H�2_ތ���QӖ��l[a��m��S��U㯏����Z�SN �1f��<Z��6�'E�o������6T�l�3W@�;1W��-.��͝*x	_=#(u��s���/��Q��o"����Y���E�0'���S����*$hW0�C�52t���A��ڔ��\�^=!6O��ߣ����GeNyz�}1���$�A9ԥ(�~
�!Kq��e��)f~�˱�ys��XT>�gS�c쨣cb57؊���q���Pʍ3@�#�z^7Sj#4ܫ#;�&#�u�a���y�����X��<�8�B��X��p͑ߖ͘��7^~���wd��C�s��`�����Rq������K�4O>b����ܹʝ'4K�h��p`M�=�]S�4�&��0>Eni�`�)e��uc>1�܄(S��ܞ�M����D@����Mmj�����n=*"u�C����.�gq�=f81Q�V搝6�r�*���џ���[��C$�2�&��.�G5��^~�ʣ�k˰�]��|�ZT���2��wx��"��4�]g"$�>�`Y 
�ۺ܍h{=C��
O�$�,�J���^�ϩ�O��|B3WD_%E��2ƫ�J	�X~��L���t��چ��p6"
���-$A	Y�����I}9�W	�^H�:��3K�0���I{�2)��z��k���>2�S^&9��1q;������k)�z�v�t Ϣ7%jq��I�D�JT;�p�V"U١���L[~��������֔� �c���޷8��)�w-�����b�:���.Ɛ��龤y?ϪS�O���oɓ!h-������u2z�.1��9�'\�oe���[�\�id�B�O4�?d�����Dq���yb�r�pxV4���R��r9�M֔]"�ۜ� ���Y��N�;Y*�>��?om�|�����SP/=�ة�*�h�����s��\u�2 �@����3��;N�Lh����=w;�z~��	O�c���8m����@*Aդ�������)sy���$d���6u�"C�0������	thp)���W�%D�0bSr|���qAf���I82?.K/q��� ��pe
���9��/4vexz��R��Ե���[v���>?>w�W[�6%�F��y��`@[V��)�.I@l��i�<I�V�A
rn-)U�O ��?�㊔�����ZԌhVQ�k�P���g�s2����q��~@�Ĩ�3`�Bs�K����$������P�$��?��"��
=��3�#BM�}���[9�b���ݿ�%u�T�h5Ȳ�����5���CK;����o]�q�,�f`�?&�O�B�JWoU�'��[�c�\7������M��k����H�5�*O�-VBЛ31����ԫ��o�`/���W:��>��nO��(X���MKR]�GhI���2ׄ��"��KK�ȣ��CWE�EIN�e�>���1�'���b?�B�A�<3�;�}�@e�o�W�zdB&@}��G����j�ҭ4�s7��i�)�֕�Q�_��*�z$�\�ay˳Ŧ�z�N�hr�G��w?
WaA������0ג�
b�8mh�gs��� ��k߬���P�bVr-.s��|�@iI��T:��F�
	����x��-�(?HI]���:�5[w��'7��v��Dܐ�VxF�z01|c3�Q�2Q��G��	��[&6pK�H��	jR|٘��-�LZb�nG��Y�X�{}KM�}[�ݕ���P�,b��8ǎ��"C��]A���Y3����b��\AB�`�4�F���6a�C�>�q� A���mf��+�W�۾�se�@k�J.�0�`�ә��_��g۶�b�����JTDYA-E�E/�5�>)H�f���"yE)�6��p
��A��ؼ��k�p��lviy7�/W��2_��ߐRH	d4vI����ʒi��p��bF�v�DH^������)��{�a>��}![��w���*m�݁6{	Q�Z=վ_�\]��X(Z{��;��ԲF(�y<���uR>��u ��j��M�6���S)Ҏ�{a����{a�Z�'e~���t'���ϐN�Z�*�('���~8���E&|r����V��Q�9v�Q���&����?�r����=�H�Y���4��F"$��s�Tɢ ��n{G�RJ<B��j��P?�O]�:wA�pOE�i�lᜌX����㦑�wᾪ^V�>;�qZ0�09�bV��I��Q�G�?�l�8�uJ&րG뗕�h��_�����*���K� ��%E��r���m/���*��Go�{�2��M-[��t����R1�P��4��o��-x/O�NQ��P{k��ٲ���|�ڈP���#bU�/尵t��6=߈^���09�����`ޢ! b���d١�79?MF=�c�hj��KPa!��A��ي���x ��l��Q����ƥ���E+R��'���̅4�bo�	��o�"P�%��2N*
\�����i���W�Xo�����$i�%iw �:��@�u9Nz����i�p��;/���Դn�q�ڲ�?�A7,�G��a���d�p�k���26(��V��X"Щ�ԌؤH$QDm�K�$��������%~ȕ�ɔ1%y��	�&��[Rs�c�6�V�1[�iF���R-mQ!Tl��_�Nd�;�š� J#�E��5��3<�:�d�\T`It4?*��녴���1���@�Zms���;��Pm*��֡�F$���P�.���#�7�'�	�6�؋���Q�]y6q�Ew���t&�FJ��x����u�;������p���`����
xW��ָ�V�b6�z=�?�(S�8by��A'�P�bQ��?�&����X1�D]�N���;�,�s��w�޵X�lg��4�ʑ�$8K�9o�b�XMNq�]��!��t�KD(;�I�dY{�7 ���P�8(�S�{vׅ���&�j}y��6_$ޖ��O���$#�e��Y�K�P�b��/2�R|�DԐA��ߖ�mT��˹�6��F���D
�,�c��!��M�N .Pi}w�n1�d��v�4뮟�1����ϭ?�ˣ����/��U5�ƾ���l$a�fk�z��E2"�>��ou�����1/�hȣ���S��@e��?-��->��v"�V��8,Q»��[�}�:j�����8��k�W3/<%j3�xb���r���Q`�\���#l��sTP���#�g�<P+ʧ��@�Q������'�!��<��Af<���eɿ�驹_/6r�k�lL�߶��?�����q�٣'�AI�1�xA&wh��Q.w�ӕ��0a��H���F�0�oJ/��4�i�k
�l�C-Ҏ�^M"2o�,[��H�P_�'��ݖ�dby��+�x�M�
��I0��][�Mρ���K�X��c�*#׫�&8������A�Z�����!�~=��x�f�t��v�*���mT�nIix�E�����"&	yܕ���8�):����)C�;)Ơ���en�����j�Ud�%
\tM�[%3�~-�{�j�lcdW�S��K�J^�a7�����6fa���̑�L	ႁaP� K�De����r΋�aN�t%�&>���@�����P.�W��}wϬ;��Bh3�N �����{�����-_$�N�ak�������;O�G��$�|}h"� �g�S���pE!�d��J+�����X��Q�8A)�X��|���<���nf�U@CO�f�n�O�:y���3�G�����=2�L��N��#8�	�l�H�5���~/YK%k��y#cM�i���o�}aV#��z�sƆ_�G��^��Ii`?-�&���{z�\%PC�/fU��e��܋L�a��v�*��vW5Y4!¥u��vďQk��}���,�򎌌ߢy 6(������лA/F�F���s;�u.y�����)G����c�4���iH��0��CB1x�m��%�[����E�K�y����^���ֹp��cD�:b��),&�o ��z���>��G�:`S�U���WT:�aʙ0�C��Qe2P�h�����cTh��=`\�M���/0%��)[,n��8��ι<MBO囄���ə)�d���z��%�Hƅ�)����U�h;F����^�5jg�W11�_H�=̕>�p#X�0f$Ɠ +��#n���'ġ�	��7�A��iHe@�w������;$?vB}.x.�oD�f�?�<���ӄ�3�3��
���\JO�ErP��hG����, 5�h�f��d~��T� �,H{�z�d�g�����`��A^�'�>���L�$����@ǥG�X�>�f������'�4�����:ԫ�"��/��Wo��f1	��T(�FG��ƭ�r�^���P^�S�WԜ��O^��r�
�����CYV��_�=��~kş(�D��'n��*�_�փ��r��X��>gЭ]b��8V���0$'�Pm�Y�����@V{�U� g��x�b�w�a����c�
�@�R�O�\��
H�R����H������5�j�#
VR�C´��9#����������9%'VY"p�)�]�pw���Ry�w�Y�+�U���n(]���N(�~ݜ�e��n4���ւ;و$����:��/I����rF���#i�c���»���R��t�b\"[�lr���=�����ǀ�7�0E��2^w8�]r �s-`}��co����Qזp��2A(h�.�d"2n,�R[��\Q\�jhz
G7ak�nC�D1.�ˈ�$3�%��;uV�΂��?��Z�8'ͨ�z��k��9_�g�h �2H��pM޽����0i�li�ࡁ�N�+��ô��x��_8#8�[|P\Mu�Ū���6\���D�醙���=���A��U���|�"�;���"�Sma�}5A@@L��.�T�R��|��^� ��2w%�z�z���@�H���k���Z��G)o��}���:`�b'Y�A�2I�!Pv��*E%��GsI�[��ES/H�����*�gs���7)�=T+�M��4�w��
�}�_Nlj>�a�(��8���cy�[�g0�d��g�	�E0X`���!�w��ծ�� A4ξ�k�Ų�
�� ��T�h5ϷXT����4��%�I�Q����I��*!��>�v�e�E��m�Yp
C�L�3�x8�7���!f.��u4��[�%ƺ�w����H\V}�΍�C<'��7�����롨��4Z&[YBm��S�i�g����������Ŋjl��cF���ki��*}��y׸�e�B�����۴����W/�h�@��8��e��7�~J�ߧY�āJ�?Cຸ�l_F[���u��u!-��Kqz��qoX����Uv�T=�X�s�<�����"�E�� �H����:��N4�$�	���3<ȡ�Ai�G?�*���ϼ�J�@e��r����T�4*�ZqB�
�_h�L�����a�0Co�S*�XV ����'�6?���_�2�5�ѵ_NH��$&��x���5,?�O�TX�Q3dQ�� �~[.�� ��͖�aV%8�W�;
�����/�0���k3���Eф�a����B�@�%�C`���dqcKY.*�� 9���¶�C�=��ӈ�j��\�p��s�G����C�n��h�0�EB
ߣ3�Z��)�/F�&�	�3�� ������2l���-p@��N�D��(�Q$u���,h�aq���Y�0�GK��	��K[yba>4D�?�`�:�/��8�9+bt�Z%��#�Þg�m�������`+ޠ*�so�Ѐl�'�X�O`v�1%5��D�����Cu4�<`��͋�1�U?�S[$�����A����563�k"�q�����/�������f/�at�9#��^��(�T�8v�ܗ��Ŵ��u<�=W��2F�]���Ė��:���{�{鼙*Mc����c��a0[K����d˺9����)8'�Ɍ�[�����1�q�5zЫ)Bk�˫wI��W��y�Q�o�u��Z�-ƙ�y��6soȉ(�����ȓJ�m�)D,��$,a[�7m��mo��(�\�1�l�s��a�'���9D��#�>#�'���z/z�����X�(X.J���y���MҊ8(F�*%t� O�8��fR���%�q:ķ4D��B?�]���-���	��A�1bDi�)_�>1��Eʖ�ٸI�U��x���S�_�M�WK���)�Ѱi�ř���y��BS�����2$"��]��@N7�?����.���B�,��L�4�zP&%o�F�A��,�m7��]3�Zؓۨ؊`�Wx,�����Kdmoz���#p_���!V^h�v�1]ݚpENj��s�{�q�q��L�8���b��l���K�`��������<�XЪP�9��h�=�=pm̝I4` 
�8~�7����I�#.7�'̑�x�x�SU]�cp	�\����V�!����ƣǻ�YT@r��;6�0�q�/�nS~���mGT�V���޳6���;V�����͕4L�-ӗ����z%��>E%5Q���H^G�ޅ�����\d�w щ�f̾�Zx}���/��G�UܿA23ddW����z[��ě��`�R8��Q8��韨���*��&���(�3?4��Y�.�At��jn����6�8\Zt<I��ީ+�d�4�6��e���/'F��+��^%��ծ^E���*G�[�7�!w�����WM�<.̎,C����)��D����柋�t@w}#�,�)�u�f
�V���JD.D7�w���l�ʳ��Qȓ�RI(/�ݬ�X�C���;�>���xh%w�l�9�J���!Dm-��۽b2��=/�Z
h��k�;�[~�lE�I�f���x4�I�A4te,A�{q�{1ϳ�_�zn�����ZZ�z�pqĦ�ru����"n�(sZ��M<Dw��C(jVZ�� �&9��|���٤�^fQ�ǀUOo�m�Z;��d0���z�`Z�d!p�7$��-��W����x�-,�B� �+j��G�rRy�����nEwE�]��E�U(�Q�VY��;驓��F���m���ة؎�TC�
s���R���5YO�Y���Q�A�y��J�9D�Z+IA�e�t�2Y9��s�2�[��gUv�Vmˤ��Tע����랝�C��R�;D"�ۈ�
�.�B��D�.�B>m�N��{�|�5��լY��;���$�Y���!��&cI+�H�FZ�s���m�:�>�� L Ե�ݜ�f���Kǅ_�8ъ������p'T}�pa�*'��8g�A�'KʊDU�1I�$z�����[��h��.s����O�w�r1���� �ݏ�'+�|}8��o��çz/Zp̮._=z��� ���]֛�ƹ�4x��Df?�W��1��y8�`v%D&G���/%?���/��x�2��MyG�"��_O�L�%�����ڴ�$G\9���p�Q4��A>Y����H� �D�*<Hǳ'�2d��	h�>so��+ۈ]��%IC��ޠ��`^܅����-��,��w�"��'*By�_�.^\��l]��� �h���Bˋ�	�R�J$�^б���!��ïƟ��p8�YAރ�0X<o�o�W�#�,v�I7o�{쮟L���W"HK�j!H�I�/��.]���tpB����^��P߮3JI[���r��J�;��^Լ�!�c��� r�L$:��Wͽ�?$�N�,FB|2~0�N˫bM��^H8+D��BQ���3S�pO�Y?�t�c��H�>��Q�]V��nJ,4��3���#$g���\�w*������a��&r��'���7]	����{T(� "O'4D�mЪ�#5�M���͕s6�HI:A�+?Ilh���Y
0d���7Fc}�i�)��D���` ��C�Ck�St�bR���غ��pJ�B�LX����no�)c���#�5̍��<	�����	zv�=2Vy-44�ML[����%8J������t��N5������mI2 �doz����4����чbhT_o\Ȣ��E;yPxӸc���禗��K��0�C�8��4s�B΢��d}F��k")�D{�>Ϻ�V�ˇ�"�=v�Z�nI4=5�͈�ѷ�H�����$�M6�9���f�b���&ec��T��#0x�wo �-.�Z����6R$m�����瑟����S���u���gB�sL�4�o����h��g�r�X�$,��i�j0�%��}\wz)�=���݆ꍼ��L�-�FlB�����f�G�ৈ �m�#1ۀ��"�q^���Z4V�z��ra��h�`pM�,��v@x"r6RiW6�MA�
����>tu-ͱF�#?��u\����ӛLD�:�r}�.n0�j��m�ᰂ4h�=��a�{;�S2����0gy+`-:���$��#��!���hQ�)���?��C�5�\��F����~>!B0�-���7U䬍Z{�j�p�dq{�-�o�8�BnQ@��(�>�a�YbC��L��N�eɚ�G9~&8�`���C��k Tr��i{���E��0�o�*`�v�HQM�
�
�L�i��T��2�ۚEG����.��^�n.bz������iC�¬mo�u:pں{���zH���ǣ�FSoG��i&��l%����N]�= 6��_*$��v���;�n�@�MÖ�L7�:Cc����z�{+��3xb��q�S��E?5'3�����Q��
@O�T8�	L}��oR]�-���]g֒��Լ����i[����B�2r`�ʊ򗋵6�r��S	s�ؚK��H��\�ݲ�1%=2SV����l�����d��E)�ԛ���@[����L�Ꞥ��J�/�*2��g�޺G�U����f>#��>�n)�02px4��Z���#�5��[�Xn�Haiz��"�~�Hp k�JbrcC��=:�) �>�	4�.h�s��Y�U�崞Y8�%����ϋ��ɏ���>�	�������q8��^�.;
�ܚ��V��˽7$��O����&�oÓ�}��� 1*�3&&�!q�g�皍n���l�w�ר��oJ�����q��4m��ۆ��С!QE���y_�Y�S{M��(�����ڿ�4�������1��T��^�>���{\Q)�sBW"�rj�搚���h�M8x�C�9�ߥѸ�߾m7茗�jN��������\7����"e����R���qG��ї�9����k�t��!n�����|��49�J&C�ST@t�(JJ{������u=PA]�[�|Z.:(�8�!:A�:o5���"�H��쳮(o_�;�i��9*c#U��:���,)ӚOHUh᳤bx��+���-!J/���ԛ�]!I��+WBJa�٘��m��R�Y��5�^Ͽk|1�L�� ��De�E��.�Ɗb��VD+�nZ�\ǡ��z�ɩ���~��h����nL�2�ܰ]�T�� Hz��؛��x�*rÖR
�����l�eT���k:^�*@�&7����`�)s�h?Ξ�ԯ��Yh2֌�4.8��X���u�#mq�W�}c�ߤ�}AbV`#ꑅ�9���.�A�c���9��s'�7����aU� 3���>*����J}�(C�3�L��)+�s۱'���Py�}�0�W��剘/W�a@"<���$��E��s��꺉��M:3�5��7���1� W-w��G��rh�H��@�Wce:��t��	%u[M˪�hw*�N�bvo��e;v)�#̐d�#�A)J�vq7L�y}0��d�r���k�=���wS=���D���U�p�����䐹In0gzMI���
F�Ji�;6��		�b�!�U`����0�y���;��)X���`r��Y?
Rv4K�DÚ�ֲ���.%Q���er|<���.��p����ƣ=��f�T��H�v�����i�\?�.cM�5V1�X��G�ʱ��/Y!�]8�F��u������D-�[�x��� �F+4���nij獂�{�
�R���w��rIlX�M�%6�\.�8�D�4���)�cɈ?U���QP�B~X9@�Rh������*��On�}VB��_�es�p�V\	���jGQ�}d�$��sb��+H��ù�����L����m�b`�]��C
��Чt��tXq?�7nM���L��O�%�����cm{���M���if�?�s=���@I^{j�hra��S����'��$�Tv/�de^�*X\�S��g�t�n8��g���>Tb�mf�l�18�'���r"!�s���"J�	�l�5�w`�`"��
-����c�>�2�t�~ja�i5��h�U����@V��d�R�%��̴>�ؔ4 u4���I�^���(�\�9�ժM�e9�f�߾���(��a!ս�1��4�}0磽�����L8$�d�h���[9���t I�[mDŋX_��O;�S�2|G�G��/Sˮ��-S���%bnkX1��T�c�gNU�@���i1U�1���to� ���i2y0�����ݎM�$i��e�!U
��ԓ��9�X��h�!2Ӊ��]��r���>��E���0-G�*A�Մ	7�h��m���?
�DT(�~�n�����
o/�
�ɩi�TwAs�y��h����ZB&�K�X"�n��H~R4���������&M���.��dZC�I�꾛�B�����jC�۹o:��΢7����]9�C��D&!C��(L�E�"�ߓgD2��+��ô }�m���X�2��ũ���=ޗl�.Xrf����J�� 
"�6+D���$�}���%'GM[q�n��.x���4'r��e7EQ)��x��iujX�g�~Z]�W� ��X�j'7�]�2��G÷�Z�]�8F�?���2E��a.`��5
�p��W�bX-q׌r3�.�[,)��(.�h��\N@��-8 kv����Oy�F���R�iT�箜��i�������%x|�ҧ��%Fk�ءK7&	�O�Y����Á/_RB��Wد��>-���|���^����3X�D~d��J���N��4��)�Y�۵�F�^�$[�u�J���|*�^�c:UEV*mQ�Vz�?�����f�DͿ4���Vw���U�/��w"��X��$:�
ك0�ZGt�!(��`��Ɩ �ﮊ.V�l_���r�
3&�h2g�}B�|���:V�*d��p�?�\}m]�'�}T{�I��v'�,Qq�tU�3�H@5���w9"d���� E��8M>�K�W��Fjf����my��`�7'��:�yn0�>����<�xB3"f���餇���t짓p�
��#Q��ϻ��'��v:�"�":g9>N�801��D��,�CV����2! Ni�K��f	w��(ϓ=�ϬW�'
����,fQ%�r�r+�$n����Y"Qаਟa�HC�٣�Wٝ���UR��s��"q��!p�h����Oت�mM�&�jz�+wKG�.�]��*�F3dJwP�����W�����Xl>
1� ����&�A=\�=M�	��9֥|T�7��?�#��ئXP�LUĒ�"���8x?�_��^�3Ï�o�����SxV0��\	�"�˔�G��	�̞�4�u��A�������z%����z���p2��v�0��|gƮ�bR�����Ub�!#u�	��]:4��P �*�2H��F=o�x/�����
����sUT�ov~@�ݏ�f}t�審8;�:=���H_1.'�s���hZk8�A���e.0=AK�,`o�ַ�0O�L��Aa�&<I�O=�Dq�/�w��r���3 �����3�{&3O\�o�.��I�ը�.�������3qq�H;�}붓G��j����@�q������dO#.�u���w����ӵ�R���`!* w:�Rچg�h��:�����E�����em*(��4}ي�8X�GF�<n�U��լn�j7[�k�����˖S�!;��d��k`�w�]�9�i�/:VQ3j�������w����z�d���7T-z�,��X-�w%|����󄔿���R����)�n��t���Q 3�)r����1�� ���C�c�7��<�i�տgv0"�˚�~܂�6��VT��%�C])�8NX�����Dm��ڇ}y��N���d��b��O'��d*�L��O�.$]��f���N��yd��	�$y}x5�!�`b�z�j�2�� ���a�(t�����1�~;�kkj~;y��Iq�l���>�3�R��m�*��Y}�6+�b���3�܋�"����A��� �*��'hV�؊˵��/�t�4���,{�ęR� oL�6�'	��m�K��Rz���t:S<{��<ɠ�p�t�@q?���g�nȧ=��e�E�T,��&�&���^�����o�#锤��e��Ph4����s���g�q�7�Ե���T�9���l2�D��Z׹�4�>j`���W鶔���e9&\��tai"��-�L�s�)����}J�E�Ϗwpx���|`ˠ��{�`:�J�sl�=׾�p�yW��s'f��Y��X8�l��p�O�8Bf�3�	�`2L�"O��I��c��ns�+KyD���;��Ą-� 8�*��Eb���m���	ؾBړp�T�+�o�����P�����<�O9G�� ~�)�AV��V����ˑ��x�����pP������b����А&�T[�"��@�l�&+��`m���c��Y�l�~榃��=s�_�b8͐�e�,+�D]���[����M�]���E��~A�D��G�Y� �3�IܺK�:M�\tC��+��z��ؕנ�N�a�is��m��&�KM�����D���e�m
�݌'���2ȟ_���U'�'�ʞ=����G5��V����u+�4Z�`A��کM��Ե�s^������DIt�Υ*l��jJ�U��؞��-��iE�H������r�bj�l٫��\�
:uIV^��U]� �k	��?�FG��j��VW>��!�[G`&'�d޿ER��C�7�8m��/��e���W��u-�x�j��U���p2�8O4$l�kx�ˬ�\���ݷ�/� ��΢a	
�O&n�����R�(�5��̂z�,�f5t4��7���A旎�����Fύ&��
j3%�����T�b��K3D���:���T�$`rZ׻-�IEu��U�3�h�?�>�\��"O:�D��ޝ�>?	��5�~���K���>�q��_y[�A�>� �����F�s�z9�r�&��ځ�����)|A�<،ra�����ژ]����0���]N�Ʒn�])`�k"�����`��ƼAoHLq�$%�Ȥ[����"���e�1h��U'P�gh����N��a^gY3��3X��S�]��(c��E��,�� шr�˴�}"�N��F�W�HSEd�8{��H}�(�� ������X\����ۖ-��H�r���|9x�i�8V���r�N"��z0���(�N�M�, �LŅT�CC"�Lq�4�����"���G��!�=����p�4���7:���e�%l�h�Ƿ4[努c⣘L����T$VBF-M�he���C*(�\�D_)Oʸ�J��[N�~-64'�:X�A��l|�=pv��lo)��G*9 4�r��a~�!�Ӊc�*����3EEN`*nk��5<�_�W���T�b���?�:9�9m��ݑk�b��PT�,��D�j�i*܀g�N�+~@TC�ǒ��������������~`�B@����U�q˻�HO}�55A�x��&(��L�k�ۍ���zȕY��X�ڑ��b]��7�˘K?�`��:�{9\�(B�I+zy	^�N���^0��0��X]�okb�bd�t�6jϑ���vKV[p��ҷ:�璙9�+����7��'���_l�}���60��X<:<��Bb�.m�*
��<C�D�� `бD
�O�{,��d�Ƨ ~�S��R ��j�t5�h,���Ĥ���%�c,�TTɖa�,���5���V�^6Z���7⺍��ٯ3n|�ʒ�WB�� ��$~��?�i�'�b�(�ݪZ[ͭ!�ڛa��{�;��ښ?}y���$ZɁ:�Tzҫ�X���{r�d�Z�kM|t�|�4�䧭eTq-�K���,�,���hER�%4����0��ף�  �˨��
����ҫ�I�Cb���P2C�U)��н���:��|?wZ�N�x�:CwY�r�oi�-��+*oY��P׀tv��W�M�E�x��?��G�Ǎ3;v����ς,���?Ys�{��I�B<,��JJ}k�R �;���-��N2�i��Y�#��`��}
��+S��u�4Y���TZ�}L�}|
_xѶM4��C1}uE�a��H_�H�K�0 �!�F�n(i�ߕ)��m�R�G��WYM��޷c_jG�Z�"w��m��L"�	B5t�J�0�"r������&D�0c��j�� m�x'f,GP�&y��%[�=z�z촓�:�Lf<u�ﾤ��3�8�k�쌽/<Lj����� ��$W�6:�=�Y��n�6���e�ag�y+��lx�f��/����H�	ס=����)�����&�_L�������$SO+�^m�bLc�w��&��I��=4s�D@Ԣ�s/��̈��5��:;��%���L��ᗵn�����J���"�&j��]F~ϟ;D�H��[3
2x]��z�.�6�$�=��UjK����Ө_���P~x�*���'/x@��u`�>c�߲./u�S+0�#+�=��t��m��p�������Y�$���[�q�:���X��FN�֧��D�"sV� ��ߟ� �?8�fIU�0�2O��|�o:?H=�VM�2M�榦��5i�K%��߶J'�T'l2�j��t� �nZ�O�"�n��G7�A���
g����#D�)R&������hL�b�mlQ�� ޱ��Aߓ�ָ��(�[��<<>~�]��ʷ�k\��+4h��#��C'���O�I�B�ȱU�wŉ�;��IzI��qvjԡ�> j�����(%*��%:M@S��F��>�(��K�3�!��o}>�#�-̵O��/U8�w$����g�S��g��d�T���|?7�n���E<�@PI�f�e�/Mj9�Aǲ�V��d>(��M"��Y�JR�W�yN�ٞ��z�K��"�#�*����:�w��2_���0���I,�Z�FW�����S��⏒a(F��<��o!��5�y�/x�`k�"r�X7ot0���G���C�ysゐfd�7�]k)�S��6L�(�Ajh���,o=Yp���C� �0�hrL3��bd?L�<��5��;~�m�o���$�����t��|e��.��#�v^F�w����z�$��! �
n�Ɵ���z� ���Ҵ���3=�(3`�Nm�L��
�a9[�F|�P��qG�L?�=T{����Zr����`�����_`_���l�g;�U�ǝ'�P�],)��\i&�"��F�uʅ���V��>����zy��\C�P����(n���}������!83$ѱ�|6�[�"���g�-�m�x!����"�`�G�� M������q{4f���q��'T�)k���Ƕ�Di�MF���l-sv�JLm�zQW�)�㖺Ӏ�qYO��'Y��FK��W��7� �?`�]��`8;M��i�R�V��Vu���ì��i����R2��`[��,�r��V{	!�?��c��WC���7 x#�9W:��٧�KW�F����i��<���;�$����V�:��T�4$�4���3����b+�;W���z�bg� �.v�`�q����7��ZYɻ��v�V�g�I�g�&���N�A��������.�1a��{� ֞k�T��v�(��/���$���� ��C��w�x� ������;(�䋱Ay#��\7)��va������K����9����Ê�(����[�k��u-�!O��~R�K�0o���=� K��xʂ�����*||3Jg�_�H��Af�3�»b�����T�k�ޠ�	�v���J�ݦf@���|�}�Y`d�R��w`�@E��~���d̋G�M5ç�3��,R��qDM��B��!��u���H<͖��М�l\ӓr��)�_�f�	���9�T0ƃ!�J_哬YS��6�k���sR@�Uoh 3^=��X�L� ç�O�i�C��U�s?F��+����e��s�}�=s�U]�Ų[�u#	Χԁ^&���0)�s�����7�k�~��8n�-@��x �v�ƹ��w\�g�����lZ^���|w�O�)��Ar��!ch,rB��Z�C
7�6n#�n�'	��˯j3xhz�fҳ��USn�l,�H�5�p��;��HV.ފT��\�����6`�U^�<�!�z-���=�:���K��2�Sr������W�6�g�NX-��'H�H<E���D=�pbAK
��N�sJ\R���"x��'���U��K�#���0��'Ta�H�):x�����Rкx׳sU@�ȹ0g5�3E���E8��(?'���b~t��0��63OF��NX@?���g=�
!�n���ԐE�=�?��!����iqXyՐH|Y,:�&�%�FG�y8;�I�J,�a[�Ǌ{�dI3*���/>��2g�W�>$3g��'é�ն؏��W2}�,m��APX��@�mƶ�n�2���aB?��&9}��Y5=M��ڛ9�R���{�.����&we�Z�T�^��E�:�h:@��%�J��Ϲy1c�Ѭ����.	��:����&1<��Y�ޞOfS�~�U�Pj�q���veO�N���x�8���;�9��!�x����,&V��!o��(�K�+���T����p����`�?Qj2�&�b
�Kb�>��R��4�Q9q�kΟN�����x���E�)v��P���y��5|�� ���g����vR��=F���|�E$���7 g�l4��M��tn��[[ege6N�>�kDe�����Ώ���i��n��N�`:y%���ZFE��<�	ǝ}�e�v�b�� _r\͋�|:Q<�X��I��L�}~���K/#��k��Sٸo��]Эg�k�[�2YTj���qǥi[���5���� AHؚ鿝�d'�����-���+�����v�}�l���mL�Bv~�^����b�S�:�I����IЦp�_[X��i����U!���{A*��ڼ<�~ɖ����P�-�B�97��%%ц����ǹ]4�)s�8��t��� �����&�Mk�M�*lW?_m;:4T+ltJ�6ċ�d�UM���{�\E�8�]����	|���q/�,Š��6�/o�k�1R����
��h�kq�x;릩hҙ��<�m�*�����+E��a2#K�"`꼥\������e���RtW�4��U����T=&��0��8�5��u�~QN��H��#32���d��=�d���S��U⋔��cTə#9�!�i��腝9Q$��|>����2�B!�6R��3N�����P�	�v�$����<�4�A_y3�{:������^��`b�C��)m�J�w�J���*I�"�11���=�ڵA-����ˀ:\d� �����R���U�� �%�-�/���k܃�E�C$��I/��r�#�8��?����X5k��D?B�@���-��hcϡi��B�B����bb_>����xn<8b�("���Ӥ=�o���V�m@^`s��c%:ٌC�qVy���FlŢ��)	3[�l��\BT�g�&��hZի�5�v%y�)O6}Б`�'�����C��йR��!\���f��$UHZ	x�@o�����aBQ0��e�FN%#2!��U�l��_(�YW8KA v1(�׾iX�6^=*l>A-�[�gq��t^k���%[��+��y>�LD�N��ի|]�c���ubOIa��G9��	�.��R�m�Z�װ��쐦r��*�|�l�H���~x����0���&�Q�m3��Ħ�,|���j -�kGu��rn��	5v�)���hG
4�Z)�{�a�K�x���<���/�A���%Ķ� IfX�ف���� ���bã���B��:�­��G�z��e���v˰���]��|��&���'���sL*�����w�\+�������v���h�Ҹ�e\�"V���у���.ri���1Jx'v��9�T7��8_���F-�T�N�#��s��R�����kD�$'�Ke!2��dn����ָ�kV����Y���(:�+al�q��� )*qϥ�p�������6U�pĊ2��&���a�4�����u���
cU(�2���)=��B���~UY7��wa���m �I'�V��5�����Ü$N��l:����| U�EϨ�u�`ڟ�|M����N�`эFO�x��~�>$�He�:�w>:�M>�u�&]�Gnq�&�]�fL�C?�ͅ�5{И�-a�>�n���$�".�Rr�k)�(<�4��9�����'K��E�����	��4���h?IX
���U1)��'�η�s5Y��r�~��1ʗ�XX�,j��3<�ǭ��BQy8C��h�)IR�Q9Gk
 i;Lb;p6Tg��!���Py�~8�r2�I�¨��=	��?�'So�;5��	P;ka�7`[���;�Ĉ�͔ȋ"!@u&����H��Q�F�~��>B��g���i�%�2�KsT��K5Jv��(��Ǝj��јl�7H�u��JQ�VX��Vny�AЋ��-cX.j}�S'����ݢ�8�X;�?�	��3s)�]�L�,C 簈
�C��؊�Ny������`B'�#��PM�I�1s���ݴp�jUU���D�k��}z��?�:+z�TO��Ck ��"e~=�N�����a%yP6�b����z�x�K�a����%���"Л��8�T�G�j��S�+���DR��{��Zy>j���p	mh
.͞������%@	;���jFG���c�S����(fqWw�ߝ�O<��d&���Q���Qn�cTT�5�b�X#�H�08l�5���Z��,wF���|��K���1�D;�>e�#�~�K�C��u�Wu�]�pN��ת����iԙN9�3�}��g?�a��[�F�P�ZTD�_�˞�Z��t$��Pm{NX���+���R/�T�V�J��V�����w#{?!}��*'�ڵJ2��П��b� ?�Ij&�;P�Vy��]�9pI�s[�ٿ�׃����Lj���k<�S��5����N�8����1�rý��/�}%��=������k^����퀂���֐���E��V�$t�������Շ~��b"A׃����$Z~jTLWa%��'7�7:����#Ku[���Ց�H���"b5DM���`P�/JUϻ��q5�e�'��ϖ�ܰ�u>ݖv>�gF���7fF����d�h;�e�1�#��\w���ͭm�����E44W�I���x��9��"YID�#��|�<������u���Bo�:ę9n����v�[�`�5��B82�Qw >�����H����P������Zv�,Iv�Q䗎�� ��]�9�1�aR_��k������]�nt��b�F7�wP6�lM��> tF�6��0�-\pNz�1~{�%���vt޹��׷N^�Z��#������5�t-\~��"�2Ϻ_�Y*q<;��x	�*7�����
��Ay������gl,�g/�܆v��7kkM�HX3��?$�����a�D^�&@��"�)i��Y�0Ȗ ��Z;���^#,��J��Y�h(ز㫂n�?m�(z\uU����}�(�����Ul�+��@q��q��n���g�Γ6�Ӡ>蟾����B�]�[˹����Pc��?�w�����$�r@b&�7{����Am6Ro죤[cq�>�_R���V�$���W*�z��;��END�2��8������f�tF�A�����,�dB mP�G�}ۣӄڥ��-jy?�Hbs�T��`Y�c�KF~�B��)y�El�`nL��´ ��jT�*��Z��r�We,���@�P1 �>Tx �;��8o�Z#i�fS{Hg�^��<Պ^�V��W���"����䥞�S!_S��O�}ٛ@�G���*�����SΌ�"��XH�;�-86�E�?$�ťu���1ү��~���ځ_M�OR<A����e2E�ףiɔ�8G�m�Pv�dDu1��y�M\NzB?�2��[Q�I �1�J��z����
���.b����d8�S�����ݻ����Q�=w?hL�uaj�$~�lȂCSc� �؄ҹ��G��!b�s�Uv__�̘|^�I;G�O>�{��OV�%�0ȥ*��8L��"�B-�e�:���ZJ�14�å�e�q���/C�'� �$Qn�X,��`�:�`?�ο�	�J0N� бZ�e$p�O-4��hv��A�����hk�*�����AP������Wu;�����\�q�@�䪾6Q*���q��r`+`�$v��m͢�
��XzC	��{�-���O�A�U��緃�)-|F�U@-��4�E9�U��c�ù��o�J}�>��bnQ<�AR����g��ք��W�D0�a7�E�A�I[�a�µf��q�ߡ�h�/nx_�����7���0e�k@��_V�}�)�Z��0ǀ�rD�H��:��&)�ņc�Z/��j!�G��I��2�5�0�7m�M�6��1Xj;F��Kr�6�/�R J��!����y�Aw�7�m�W��R>�A�q�R���ӱ�Z�,�Ii���a9����Ha��1�Q���sD��*<71l�FB���'8`Rf�����|�t)�X��/�$%���&$�N��J����g��T���q@���p���TN�	��v{^7��/WG�an1r����?|�d��<sn��զ^���
�!�R��ƌ'P_�
�{4�:a��_�J��I!K��bM��J-�¬s|��Q���.��}�>CQ��k�o�a ����F���L7\(�+,�މ�Ck��@��a!Ѧ����0X��-Th��\{�~�E��]Z����[��KD)IZ���O�3+�F����]� ��q�:�X�	ki�����Ǎ���e��-M��� ��I��3u(�h������,���k
���V���Z��\���Ҽ��5��,�
�x�w��j|�����Ӭ�.�{Or���J��������	v<�Y@!)5����G��7�Scf)%9�ܢ � ��<���P\3��t�.�5O��Bϐ\�+�r�[Á߿�ݦ�I�C�~�V_��o\X��;yk��ߧ�g������-ՎgL0�,��|�rL����	&�#8�$O��Q���f�����F�Ŝ��w$��w��(z�ӠMҿ�1s�-)�iڱ��؃1�/^���(/ƻ7��[�4��)r�o4�܇ӄt%@Μ/��tQ��o�T�HN�&|.��N�փ[˜���Z�0�>�����ߔ�T�WTܚ޻a�|嫣�*�0�W%��aW�#ZN�d�pQU��#R��{^\�Zt�P�����o�z��ֻj��ۮq�����Y��FS?���*t��Ѻ�ĵ<(E���a�6�t\e�]+��2�ې�_�2����Otwθu�.����mF�r���[�g��
����XlT�F�M��P��9� 4�����/�C��|��3@�v��Jf�KJDj�"���'�d�76j��&ϙ��@��gcVH2	��IiU���mK�9&�0��Ͽ�b<��JR�@ϑR�=;�g�����ój��}J���5�����5px	;ݯV�.��&���d����%���pvh=�}�_�d���.J2����',?��ǂ}!��9�R|�z?����f�*y� �r��9����p+�^��`�꛾Թ5�<�c>*�>dt�iMP���vO�R�N��G<z��g�JM(YT��\�oLR���U&�2
Xg�id�h�������Zv���.NçC�����KM�֮ypA�{��c��`�p�&b� *�ypQ�D�=B���ݫ�ʨ킳�?��k_�0���3\�y���U�Z���C�Zl���k�I��;S��x��l#�� j��[ӳ�R��Y1W�QNB�yq�H�9����	8/鉎�#���p��D�D���"�>K�y;��Dv���c�Ԅ�ܭ㯄��������F�+x؇�P�#=e�e�-�y���n�� ��^6O��[ǒ��.?{�[}�n�H��Χ�:�G@(����S3�r�1}.��zɆ�ŷ_ni�A�ˎ*.7k�K��R��-r�S�ً��ŃՉ�C;�w���?��y� �� ��Ǟ���:��������[��pRȈ�$te ѱ)\��b�R�r�U������t�z`�fc��F-���#P�^�����@7�V�����?#��ZO�%zTS�\Ŕ���!_���1�^�X�_4�Y�p>�h�)�D��IP���}x�X��:��u�cu��Zf���M���:��<3��8�R���p(�z�>k��O]ݵ}P�$��v��1<g!j���wkaϺ(N�����ʜ�M.�:�3Ee{W�G�񶢊��"�k�׋�7�j�͓\/Z��P}ƐDp�e�w{;��O	^m����$����r�ky�K��z���r�s�|�����b)	��m��]�|�C���,*��O��`tX8����.��>�x�A��" ���gl=d�^��U-�QJ��������C=�e�Ł�h��9>��[HJ�@�����*ZA/4�=��;�q»�T@�В��A�bجq>��?Ґ�J�{2F
�F���)��Po�߻H^���!W�L��nhl��o��`�Ն@�)�&��~��z��'�h��c; p��3�ܠ>u�p�:\q�
���D4�׫��W�_����Dɸ��7�4y��Q7S�'p,��4a����O{�4�sÒ����F�܂��߷t�+���zY��5�X&~��Tx7�<�2ŽP�Ս�G7$ե�LC{J��I� p���5�p�����ͱiNNH�����6�pۊ��8m����]A�?�t��lv���xB�,��|��#������D�#��Yd��Cj��S�����K��P�9}'�#�]_'�Y��X�(���1�]f�	�m���(~#���Pŋ����x$��B�����w���^�lsiБ����(i������m�;��5I���si`34o\�JD��za�u��^d�L;�����Z�0N=��}�^��|�M�O�,]\�N�Ɨ+;Y���yE߅�A�����3���ĭ|Dg�j6�q���}�#��E#�+\� ��H?��Z1�O?���	f��%H��r���g�B�J3�j�����~#��03n��?&�[�ʉ�t�z��?A	�^?�F�HI��_�Ng��ꯦ�;Fӗ�a��]R�i��r+B�vS��'l�����?�U�֨.��iB�c����{�3<(�t��)Br���^ب���y���9��9yVV�l..��߷>�]���-�b֛S3�3g�w3�!�#�v�c.�hG�(��v�W��Q���O@���+J�ū���"�V	��k�t�d$_xI�!֟�Ƶ�����~`��2c �����D�P�8/�����z"F�[�$�i�졖
��s%^�HR"�%��2N���ͪΖ��k��'nl_�X�x�gp�ךiW;(��ǎK;"?R!'�A$�{R��c���B����8�N��t��qWy�ٶ�����S��VZ�����SIw@U_�3��ֹ������5Ryx܍��cr��O7�ʘ^.� �1$�\Q���6,u5�d�ǔi������ゕM�r)��lT�P7J�/�Ŭ�?�U�d�Q2���N=�~�hh�;�s�C��d��jO�[�@��o�e0�r{{b�f�)G��j��ޮx�qR����f�YR�WϾE��X�n�}�H���F����c�u����\�ઍĬ��"|vݍ���V���)��E::Qj6�EI>��H3�"%Çs�Z�"��xh�S���Sj�w�--��|�l�����o}�7f������5�G�4�"4^����y�IDW��Cg[yB�
3��j�����\O-}�3�󓜸p���E�I�*��_�x�BX�����Ղ8��<���`�0y����D8#��HuF M���4��܀EI�Y��-i7�����`���ي��^���:�	�(�u;b�����a���6���f�Y���8�[�K�#�悙Z��Vd�4�a����%�K�6~�NI�_�*�jz�6�� ���.�!	4���yy��6�=aFܸ{�:�i���o԰+�S�w'�-p����'����n�_��_����������O��5BK\�O�{Ii��l�+�p?�eV��3�YW���zf !-��{8�80 ,@����k���"�� O�g�8f�)ѵ�вD����}
H�N�2q<�Y`��1D0AhS��$���͹�2A4nH��ۊ(��Bm��$�go��sm��C(ՙ���k���E)*~.6t��}�r׃'������E�m�[��˹e)����l99�� r���2�`Y�rRm\���S��f��[γD����L��Ŕ�a������/��(�e�U�e��R�G=V�F��!��`뤓$�����dν�v|4�k(	��8�s�9;�>�����t�竚)�C�(ōI$8l����PgO���w�B �ZP�9��W�3�"w�?��~k����\���g�j\Y��J��Y��]\�C���R�p���㜗���,'�\��.��U�J�ߎN����|+6�jo�gn�i��􋪹��4�6}Ie�ް0��{�K�L�?��ۦtI/�����]]�ό�I0�H��,і�?��i��40�����S�<G�*w�gm�ݓI?vmI�4�9*��L#��@�������_�!�8�a
 �w�-����ady?dN�i����0�/O�/f��f�D@�����WO������g�h?����S%�8���$,�w�:tv5���t��w������t�Q��%���AI+*�v-��H)MP�����5���%@�:���j$�U��v�`}��&�?֫~�u5�|h��4�}q>�-��ukܘ�m/�����g����gP`Ӊoαڽ����^]���3d?PQo+��c�杞I?���C��g����8M����\��%�x �VAX�v��l]��CI���{݈��g�9���b�(eJ�����
x�7��M,�D��//3 �ݶ���Z�/�M(���d�ѐ�y���	2�ާ��@ �[�����i6-lA�E���]���E;���CC1��'Z�N�r��p��: ��z�x���9,��r2m9�>m�FI��?���[2>�(ݒ{�rz���14���r�ׄԗ�&�8o�;?�tڎ	�­D�=�������Լ��9�y�q&�j0��ِ]��@��?O�=�
o���X�t�s�"/�ҡ�G�0EC�g1�;$�9A
������Pg5k�ga���
ؼ�=5�o|�@rN�}�9��Zh�6v�u�>���1%��fi.;�Xn3c��R��x�Ǚ+��/u��T� ��ʟ�F�<�T����&���Ua^]�I���s�F����*�����7�ڮ��P��a�g]��/�͊���� � | jql�[�4�)���
���B��gT��l�����4_:�*Z��TۧӇ"�t�2��a�wQ�y�Ac�E�1���9T[�0�^�ދ�_����w<���x`�F[��č��2�{�����7�ؘb������`�朠R�@���Ͽu#Öo0��B0�X��\�Y{Kx��ui�,��:ifH_�p�$��'��:�y�a�w�F�"L�;��b!���meO/1WEY��Ё��Q\^��׳�*5=ܿ�v�m�a�.��- �S���R��)����A]0Ʀ�}�hm�Dh��۫;�C;��bY�.C�`t�ø��s2���^T����4]A��$I�)��JN�,�v���x+A@�Y����xL�>�h�.NT�C�G x�%/�ɡ�Y��񽯿�Ь�B�����ƘA�����:+P�����uvXD���?g���hA�0��7��+r��������ﰠ&�����p6�`�R���i�H�@/��zZc�,�]�e�� t�·=��7ʙ젷�2Q�G0+��z"]��9��l�y�iLAz��HǗ{!�Ȏ�nW>���Q���1P�އ�v����rv�N��+���:�|ut����3��OBI�˃Љi�f��r��5�B���.V/U)�Rg��r2B�2\c?H����W�]��z������D�n+/Ӿ��@)��E�#q�����h5�y�졝t6t�o+�G_�gS�]m�pk*H�d�b����[�����]�1\)���/�[�	'��k�T�组�Ƒ$H@� 3��8Q�2�jʄ����<Tp4nd����R�,7l�$L�H�W���^Rn,=�.�N��h���6y����|Q�����8�Lq3�T���+(������ꡂ�'V�O �ݯy5M(�	3?��3�Ϡ�-���x�.M������1~7�c06�:멵�ڮ���~~��-����sk��`�Ͻ|%iWxp���F4�x�u��yU~�&��b�(�#SI.[�/5]�8�N�:��n�q���H����C���θ��W��.��Y�޼�z.�ѫ�'>����Rٕʰ�/� �G�
c�Xwg�y�D*����aC��_?��%t��b֎�C�Nru� �7�x����3����G�������bs`ہ���R�t�.��ّ��,�>�3 �,�+�U�+��w�*%�O
�����?��2RjVwG����`8s��~��w���}1�z=��N���Æ'���S]=�ǽ�����~-]��dyS`]�V�1]�tW�*�D֍�p+��g�����d�,`؃�	������+(|;=��X�~S��]�+@���|O�#�*)/��3�L��l�p�=z�.��e�J�_����v	�.4:�jr$� D%XMɈ6#��d�x`��N�k���m�ͮ q�/���q{��5m9�C- �?�G����p�L�S��s�f�mB��F=�L��I��T�~?Fq[+�gn����\=�1'@�/��k�ssw�פ� +�(���BZN�LY��0�WM;��L'zO�"�S���XJ�;�|
S|'��_H�>���F��`(�D�0���>փ�~D�
m���	�����T�ba� �}�����P)=��K��<�,�f�k�]+ � �s��,VFg��>�h�Ĺ(�t���f�]��ُ���+5��˅�&��p�![�`�{pw5�U�� �ſӋ'F����?�h1����WȖѩe	�a�$��'�pU��GDm�E�7���L�}�}`)���R��/GH��E�~�h:3�0��P�jVR�Y"����x� �L����+�&?�%DoG�H���#�}��ڽ�	�È�͵f��s:u ��sC6Ȧ���N3�gG�uz�C�J�h���VE[<��N��	�Cú��%�M�4kx�k!�
s	�>�v��Ѹ�dQ�b]���(��5Q�7�iV��m}��N�P*|ck���KƠD�>�^F���\a6&�}(�����w޿�0.J��
���{U�T�8��~��,?�2 ���&>�o/9Ʃ>!��'Lk���̱˹��q@��Ux������Dk�R�-��T��P��B!���D�{Z����kb�����ԛC)(�%EL���o4�G��&�b��Ge����b�9�oi�F�{,��Þ,F�c6E��¹���m��!d���T��9��,y�n����EA��;,[:�Y�ˏZ;�,M_]S*����hߙ�P���l��v��y##�.��ŨQ���	0�� �<�T>��0��hy��z��,���	��k�^��ġn�.�?%��7��j6��=�����ܜ"��	mV��Q���Z����+����5�їΉ~ui����nh�L*�c��CY��y����Sry�d>��.������ORE��aEJ�����'�W�h1#�����Z���d��O�7 �#T�a+�{�mT��T����j4q�z����f�S��.S\�q rj����p��0�)���'�j=A,��>�b�{���#J��3;�3�����Sq��w�ދ��]LmwY1�_��8���Ԓ+�.~^�I���<��f�d?����2�N�GxS���8CL��7�-
l���_}��UW0����X7g��Tu}u\���R�fo�10 _A�i��Ņ�=~W��{:�ύ�N�Z07�b�D��ȗ=|�d�z���M�L�14�_5�D[��qW{wUp_n`�`�xIC�w��uu~�����z�%���!-UK�s�9-��1���5+'ޯu􋣁R�&����c�����d�1DC�V�lgx<k�(]�3���	����+��#?Kک|��s��椲�F�5�;���V��B��w�s���G�*1Tq�'} ��Dt�P�C�Hu��I��n��ۈ��u�<8�y�T΍$q��K�8>���zɋ+�ѩ��SCe-��So�Z��/��-$�S�n�������}�n3���IҬ���T�~�a�c���٦qG5�o��d$��K��11�5{�3�[�) P�4'�� ;����<����Ҍ����A(K���:�}���Ԧ�*�pڰ/���z�P&WMs�{��z$Ū��o��VI'z1�Q��thn޺�l�4�c�+o6P�����~l���`ldF��֪��\������^Dh�"���״��zά��I-3�	I��v���m��:bU��kH5�Y�I�Fr�9<�
X��ؽ��nҹ��ShLk����+�b�!>�U�ǰ�*,�����a�V��Ɠ6���S��Ĩ�b��P��w&u�ު*ܥ�Y�+YB���ye�D���"y��~��/���=)�|�<�~�^���FFJ�9�`�/wܷ�~s-*c�fG<��u�?��;�q򩢤w�\��5d���W�d�jE|��GZ�3k�=4�5n �/l* ��/�7K��N��܇p��'��+��ƩF�jY�/}�袠v��� P�$��xdp�(�7��5�zIzX��൭�C*�68ͬ)~75)~�$���."F�y�|e�|ʛ�6������C���MxK�r�՛e44��T�?���/,�.�{~ry�5�Eh�t����5i=�(��΁'p�GV\X*g�g�̃�Ǚ0�Ő��5�ĝg1,�[ʜ2`�z��ECo8���e޾�)m�C�����\��ێ ���R�s	3a���<�IL?�mU��Q�z9a��*�i4�]ڮ@����k����,�o{�{6(�]����a6-Tz�+������24�ƍa��U��M&���ONbP���ї��}�i����\+u�n�M"m��E>5Z|YV`-g�]<�O3�{?$�~�J�j�R>�Jl/Z䢻i�����WX+�	��W���:^]�@q��؇���F"2��阹g�]��:��,.����؋;B� :\�fQ��e��"	>}+�Y�,M����"쀼�=,�f��~ՙ��e�@=�9(��)���8�B��*{?�4�E�m>��՚�d#�����(s��%C���WH�I\:r̺A�GvE[���7X�`�D*M���m�g��C�D�d��Gw����J2�}T�Q�	�ȣ%	V�`E��l�>غ�:�6��y���1��l(���S�^1�R���U���uz!E�m���M:$n�<��%����(�P"v�� 2��yy ]�O^С�{	����� ��h�o(�x��ZՃ-��Nݗ)�W:z��Dr��z�g���gn�]��Ϟ�0/j>Z��At���ڋ��v�2����:N��Eu�$`��)��-���12�b��6���a\��9���Rs3��-�h}C�{h/f�"J��k2�����_����<�Ӄ��8�Ĳ�������E.q�<آS0�\����15�Z���������JD__�
z��>u��pˠ_~�Y���Y�`�"�����'*�2�P�Z�ji����������UL����8n)ЂJ|1#�8�R�|����t~O��f�~Ryz�))���.p��5���A����L���9w�%�)���p��xs��#�����ByK SQO;y�R),M\ ��')�I֛��@�20� ����d��]6}<~��y4�ɓ�H	N��ʴbsz�v��Y� �G���n�
A�Ue9g@��>��"���Y��E<��V ���5�+3~l��K��O=S�2��/)�Z�<e´9@q<f�@b����-���H��3��&�6����u�6Z�:V����֭�ۗ�����{g�ԏ�%ܷ@��
m�q�5�֥;�s�d�U0�r�A�U/�<�۹�^3�jıb�TW�P�*��_���i�q~�vg�L�=���re)N �m��[b�kb�y�0���@&�H���I��${(�o]������ښ�J'˙3_�/6�zRN�{�	ڐYضW��Ϝ��*��Y�E���n������ۙ�u+*��/�e�:�p��f����4�?{�<>;up�j_5>�,~r�|��#�y�R:�6PlFu崧�6�^�2�����)H�c�w$n�葔"�θ�7�.$h�#ˎ���L���^i�	v[�	��hg�@��=�>l@���@���d��I��+%�]�k�%v�J��XVlck��DkL���[�^|�bUםދg����k��5m�\1о� ��!A�s^?[�OG��4@�%nw/"�:Cu'y�����D���R"�^>O���l��`���xK;4���Rk9ipPz���`U]#�[�x6e��g�h �S�P����bT	��I��c �݁����d�IOۤ�5AX)mW��p)�َ)`���\		 35}�t� "�3���&b"(4�U���M�T��R�V'��4wr��IU�� ��a&hؑ�n_�cK���I��q����%��O����{��k�;�e��f�[SC����\�����[/�o��u�F�EK^�`*���?6�J�O�5�������X\�ġyv�t�v�+���ӄ��sB��wXR���eR��=�����\r����*�Ig�&��L%yߟ�%�IЌ���D����J(�QV?O�� �x��H��	�|g{���5@9���bn��Zc�l��Ǧ�����-'�O�J8sBp�����}Yܾ�\{��@����q��@{R�8���L�2��\����tl��=�r>��� o���j�L��| "���{7���K��E���*i���C�N��u���� !�knܪ�ͬ��磀���e�Z�OA��B�k���I���
�oB�M�V}���!+�Rv���x˳Y��ϫ�:,c-�@&Q��,��ޞ)ih��j�G]�:�S���_x��Q|&U�lT�X�=[�\~ˠ�H;�� f#���P߻�_�ߴ��d�=R�i���a͝8*��DC]�Y��|��������U��}5�BJ6�}��ǜw�v"�O��F�)��ɷU�*3Le�L�&�E0Lμv��5���W��ͩ��;/��M_S��xw������()ÿ�����
�y���ᶚ:�bK55gw\6�+.�բ��.��ꪁ~gCp E���
XQe|A���/����v��8
���{4��c0\׵�}N&�dW��n�a_�� ,S���P)����^�յ�!��hP=r.T쀸7�].y��MWN�_�]�v'�D{z֜u���:e����Y��H_h�̄���l6��*ܱ���Tۀr���'�ڈ����1�������K��?�܁���r>��u0�%�_�'��/�c�V�A3X�����ٳ����c������p�U���f�!4��'	��5p���H�|�+��n�G��� gx7��(6#K}�Y ]�wT�|���;�d}�I�4��g�/S��!�OJ(4S��q׋�ZK_��5���K]^|���q������(���/E;eb_=�7��ަ1˔���!o�mć�"Fa{T�<�RB<�ێ��6��g��0A��_���-��%�t��%6�mys��HQ8�OfG��4�It�;uW)45�؈v��PA���f�4=֧�k�� ���k\h4@�����zjl�����J��K�����D��.����7�Ukj��LW�e�=�^���x���~�Ծ�[9<���f���T�����2F��>� �D���F��Ep�Cp(�.�]k���]��=_f{?��Q�1O��#�)�Ŷ{�=��iY�c��C6P�E���o�*��|�H��u��}��*���g��t\�юG~
r�1����R�g��7X��K��m���8p��EbK�Zne�8[9�Sjc�h��?l�:X�J�a�1�B-�\����	݅H�K�f�����rs�2��a��BΙ�lx��J�_�S�������A���K��I}U�{^X�%n9�aϿ�:��q���t����ǯV`3Y!|0H�W�Jm��٭�y���Ki��]�.�7U�����Q�A/F��:QT�F�e���K��!��O5ŌC��Cz\;�ܮF'ZZD��(��qM�@܄��3������s(wݩ�4z�'� z7/�ڍ.X�>�),j�'"fcȪ�3�^g��nG��w~ ����H�GУ>�'���� x�@����0�\�̬['�/�c�O�.r��~�H��i����A+%��s0�Af3Xŗ��&��e�����Y�,���5���A��8x��J6
@�T�͇>Z*1 cw_���X�N��1T:koC�5����N�w���{�\�����f�I�{Q�"�nh>���/`�FoHO����|.�ln�VF�R������(�?iM0����R8��c،����-?~W��Z�/ �u6�PV?�P��%Rn��K��|�ɨ:�w�Wl�ɀ�Ù��8. (�C��\�V�o��+��wI �D�A:�Z4*1��R���;����=�3�1����DH��������R�7���2���1�{��D�}wb%r�N%��2��/@I���^ngyp_C����=9��<��
��e�O"����W":�5D��I�6��AU�1�������6�'6���H�A�H}�)�pL��MQ	6"ha�ݾ�� �73��,��H�
�r���U������os74$�geL�����E~z��}���H�5HV���?�X'B�g8E�p���M2�Ԛ���[�#�c�?��V��Α���(;�~�KL��íQ����!��-�3����R87�}�m+{c���~��oR��9L���&&��U:fd�+����-��+�� b���_e�}�o��~�|�ݽ֩�j-�nO3��i!2ٚ�����d�>����q�.�H���6 �sK���ՙ5�������8�v��l��؁S�&���2�(�m|�C?�Ԁp�!$-ԟy
�c�N���z0�V����ڸy�t?1�Ҩ���ƕe$B�R��u9��$���3"QV�C��YB��+L�d��nz�X�7�#^3,�����_�X��j3o|Y^�����(����MS7FE��<&���|p�@����~��zT	⸁8VH°�7׏�+vE7$s�;mRTZ�z��h��wd��)��"����C�o�)�H`%\H�Yx�����2S�����v	� �A�+�����k�5���0q+�ҴA�VM�Ӽ�$!�Zb��eX.eb�)6#�[���W�j��A�d�n`l��	�ˊJꨖ8�|�z*O�-넥��X���D���'�t��e/U�|�lT�=�dw�-"G�0����ңi��!kw%�0T�[��bE�(}�D��a<D�8G�{���"!�z�$פ�Q��CE�hm.�##!%�2X·k �.��������O�*s�ց����� E�82a�ĎUȜ/w`m��bɰ���B�~�Ų��"y�Z-������E�ZË�^�1L�&���-y=�[��]�Fs�����wsc���><�����]��9�H��%���j	7s:�7�����2�H��)��s ��z1n�qk��æ�,�����	���e�.fMǕJ�~ V
, gTM|��8 �@Y���Ȍ�J�����te-#�V��Z+�00�&��u�RŲ�R�p)*��������).�DW!�E�7.�q���(X�l<�_{�o*�{@�x)��`�[��Rcm���L�.�n�3YTm�0��(�5�4�)ƴۍ"s/ͫ��`�|h����}C0ZN_9��.Ea|��YOv86`�W��O���T����
���<V�z6�|��t��o���fy[����!֍�D~ 8�Ʀ��YZ�QJc�!ɝ:��H�7�_�Xj�X0�F5E�h��@�ͣ��ح���#ؤ���ߜį���J~�(�UZ�=��a���������1�&������@u�|7	4=D{u�Pp�[S�_*��h��S�Ɍ;��0+P��^Յz���f�)j���$��a�B	,��6jM��룖��=�����8�gnl�Α!w����T ��y��lH2f�`�������÷U�M�N�L%=��v���,@�A-?(�&�#�*���%�̆�I&>����S�+gH�1s;�w��t�˸��.$�g�#�`�a�u�ʜjU�>N��O	5�0�O�S߰�L��4�t��=�eհ3�߃ɡ���1����sw�P���L뉛��XsΡc_����t�f��傩�`��]�>���C��=�z1�][������d?�%F<<Q	
��L��Bym��Z� �]�T����:��v/��f��I@v�z��[�@(I��%A�w+ӱ�	�F�)i���I!��JP�:'ӷ��n��
��]�-^���IJ�AdQ��!�|����P_���[��J���j7G�J-06n���B0`���tR�X@���`��;��(��/Y���6��KG�%��k��7	B��Ya 8Ϊyx�Ke*l�-_�P,�Qz��B��C�V�e���%.=os18�Ŧ��c��t��O&s�ח�뼈�cY��_= ��N[=d��6���BT�}gjm� �P�����LYɢ	a$F��j�!FS.w\12�b(�-�<��~x�Z�D��bnO{:���k�YJ s�^��^Vse�o"m0�$�����_r:����_�M��j���a���u�-B\��Y��3pǬ`w�_�ĨX���u�d��[L)^]*cJ$��]� Ѻ��tz:.�ϕR�t$j�1��3I�!���]x���u�YU��-�	����·�xӦ_���WͦK,�o�[;�����f�ەez)b�"��O���lU?�y��XFe����g���>J����g��&�40[c�NCbP.k�׺Evn�c=�d�g���Ŕ٩ؼ��'ð5	j���ԃ��5"��=ph�S�ʝ�n|�U�'JS�>sg5��.��%g�)�+�s0�wX�S�#<�T?ʿdTo6&��6��+�;����u���
��9�]��c�?�GnyP���
!�I~����-��[�~C.#��:����~,�w/�+}pu[O���T,�j3
쉜���~����V�� r��ڨ��Ϣ~&��3��/�_����1�ݥ�ӟ!���%|�ѲT�]jXx�&�����H[�������BG}����O�w'�_<�S��l��Jg�/�-բ5*�AVDI7�]N�sc<A�vj|�U���T�^��"�I�L3��_Y��U0����	�
�����Ȟ'aF���r{!&M+b�u�����f������Pd����t��{�2�O�s���3/[�͊ĳ�Ea'M���4��$"�pY��6�\-�������F��_R�H�nږ&ڔKQ���N�yX\�T�HC�=(�1�o��U�]��ʨ�x-�Vբ��F֢zZ>�����8}�C~�y�7S�:�1ۺ�A�m��O�3줿�]\ή���I��]R/6��;�LQ��wz��O7z`,{~u�RpN���������Bs	���q����XjGE�]�d3�J����R0,����A�!W�1�4�0r�/�g6� 2.�g�ۭgJ�e�9@�gU���Co��j4����檀�%�Z���4�hHZ}�!R(�3qj�з=�+)��bm��lgU��:�G���Oz;�M}�+\EO�5���@NX9AM�jR�˷�ι�9 ��ؑ²�Tr.?�+�:Tm\0�n�*�'��@�:_=W������� �]���{2��َ����C����)�*���KBa�9���Öz�՜mk�f�Z��4/ʋ�-�)�t��ME<�,��r������z.\��kʰ���n:�!��g����]�
��Jq���uq���Ă!zU�d�p�]���k��9��I����B���8�����L����cc)<%6 ��Ex��.����Y���Z���7��@X����(�w'k�%b���A��1;��w�i�<��D��A�ϟ�KOG�Ec[������}�M�^Yt`2��َ̥Y�DX`�)�y�S4Uv~�4?i��x�����<��m��"��U�J ��E�hpO2PA#T�K���ؚ�]���;X~l��v�����FH��c��M��
G��{{��󗸢��s��T��=Q(��j2#��~��wU�}�t���)�V274B�m4V��%Q��C~�*�~��~�&~�I��pΌ��y��W|�!�Ne�H�J �o�ڀ�E�e�<S2nr:Z���n�VB�.�H����I�y��u��)�DŤ^J1�����տ�e���L��Y�L7�Uڵ129,��O�"JB��;Ps����(������y	p"D+�]�4��0V�;���U�e"�9��K,f��B�Ȇ�S�B�b��DBU!��J�����W�Y�ǟ��i��ފ5�?,-{��D���ل'o�nq'�Ƀ��i�El�kx�(*�`�� \�@��P ���- �y���e�|��PA��(��<�	|?��M{�`���uI���+��&P�anf�:����Y�@����)����I+H�3X2��G�	�2�*߳�I��j����b�|x ��+[H��zز#lr=�S|�[�O��R��
�3CD�)�*�a���a�v�2;�K�"�6��`ޗ���!b�n��>�S��F����4+^�������2Z0���Y�+!�Z����R���f���/s�s)P+��y�~�m�Ti9����d� YG���L�JF\�4���0��z��0�1�^�٥M��`M���f�D*?��?��s*� z���K{7-H�زG�]/1��
�n���(�1E��D��U�z ��4 ?:�A�SwjP\�1�#C�+P۪�/ےB�u�q���(d�p��tHp��#�ê�@Zk�Z]�H�´�����-۩z"E����Ԃ�@��G�!�N�.{pJ����q����_	� �����b��M�5\"��8
%���]=:]M&��&��}���8�;C;1fЊ���%�a�L=RI�ܿ^;QL�\�p�1����Y:F���^ e�J�!�D�l�}L��ل:�mo�E՚���Z.�ɰ�}֤M �@>���!v�@E�ӏ;vW���8�â�ނ�i��~��6kR �T&�)Z6���O\GnV��;qsTڶ��6���Q�fcf��5 �|}Aa����[�a#�ӽNG�0
�5����6FF�ʥ�dưW��f��ɓ}���c7�����\�P��ߘ��%\,� 遗�����o��U�<M�H���q(�Y��~�"�I�_^?8�L���M�^�C�J��vz��r,o��w����6'ob]�}�`�П�ì;�x�
1��r�{�<(s����������*�v���BWU�iUm�!8�F�o�w�xA�o��;��4l^P��+Xu=x8z	yq�uL���n}3<�Nz�c2����=+�y�nA��R��8R�CjB�q2v�K��r�\߫�\'[=P��^�]Ө��H2h�E)�di�=.�3GrM�N�OcxT�-�'��6�]���X݉U��`�p��I�Ȕ��S5钲�ڂ�S��N��tfÊK�����~�-Y���9�AS�����0��d���u
�'�{(YN*��y����g@%�'�qGJ�+��y�疎MtP�v��h�ހ3�aP]zۗ��ev���<ޚ�z�)F�/g����w�$��E�a?�?i�Y�()��sEeA���y���6���1�K,
n�9彸�`Ǆ(G�粃-�o5�sQVj��*�k٪q��Aom��x���?�A�A���ѺT����$��W�\�nP:�VWr7���DjwW���y� ��L��]]�^�+&��8������bV�� �9��g��I�i�{�+>�8"��uIk0�ergW|��dt������V��Y��j�,J����;D,9���oP2ѡ?��*PNJ�R@��?��*�C-$�����;�M��b�$��z��JQ�0�VTDL��f�,e�<T�����_��o����R!��@q�և�B�\���#H�v)�1���U�Z�&��>M��N��Y�����Z��,%P��]$��9��
���`6�`ah�5�9������{���Сf�wX�ef�KA�y�U�<�?�da�n61��[Y�9��fbS��e�(�"��:�t��8$e�$����&��8а/���*�4Z��g��""��}#v�y���o�>�#��{ �Oi*_'���Z{wJ<��l%��wP|��z���A~�ȍ�W�4�a�WL��Rp����`<����9�0f�`[���>�H%rx���@�#we�{b�0�Dǀ�d�d2�g5�S�WrM�z�vT��w0p�뱏��B��	��CSD��e��Ռ�G)���//)T-�Зq�J���U<%�Az�H�\]�v���o_�܃P�]ztC�/&�Y�=�e��� ��B�	BA�oj��ٴ���������+���N��k2�2GH�Q���$�v��%-y��ݕ�J;�g�g��J��;r7A�w�Nb�mT���m��TkoB̨�C�4��h��Nj�k�񯧬5u1q�4��!�����!�࠙��4�6��W��Ae#6ʔ�� ��O���*9"YHI��c����E	��󘈖¨��Ӂs	K��,��$��dp.�,��5-Q� 7i㋐�9��o�d�eG7_�U0��V������V���p��p�Ę��=B(xv�)�r� ����JU�c��,���g
p�5���4�'�m��^7���q]|��7�W㧖�b��ʒ��7H$1 �'���)ƀ ����#+���.䂎��.WVNi�_197��P"
���T��\�^� MΝT�v$�|��A�ΒM�s��A[ R&��x�,A��͏(����mq����jh=��A�yFI�5�R�3P;�oʧ����� x��DxT�N㔶������|+�G�D}�	a�����izz��뽆;�R|0��Mx_��p�ݸ,0\�r��=�i����'J×$�I,�����2�Ѕ�l�ǝ�%)����}-i�����Zo�3r;5~�NX�$|���n3�o9��(�5Fg_L���y´dA1E�<4� i��g�\o&�fq�sL�����Q�M�c�`�g���GO���Zs��䏣i�����<�$��_~g�8�F�]��-��;�V�Fd�#},�˵�N`!Ge��^I�_��w���7�M�Ė�}5΄���1V޻���ak�W�<�߀8_]�v�1�I	tb[�N�Ђg"�wP��"�x��.%�M��O�aǌ��3�yoB��A Z�kq6�Hl���G�`�bx��{����#\2LO餶5���5�8����X3g�جT�t��`p5�O�L0в�H�S�'3�w�t�����|V��K�h��T��e:P�U6�q�ܺm�%��/4��V���.�Ad�b���k��f��f�l(����o�v��&7�e��/��.	���v$�}GF7�%W�/�17�d��A�u�Ұ��:%�1��<ް�������Wڐ�(@.u��pU3��ļam��1���h!�����/۴zo�9;g+���$�3�4/{RثH�XQ�@瘍�үiz+'�Zq#o�ѡ���N~��q%��>���;��լG˃���Ÿ��Z���/���D��|Z��?�p�蘟�����bF"Q~;�a"��Gmy'WL/�p��=n?sY�ޝǆX���`?u:��!XM��P����pko:�Ū��+�UMY�egmE]�ż�>�L*Sh�G�+N������6<jN�IL`���KT�<�8�ipm �rׯ���c?�ԁ����r2Hܩ��a��S�W5��.A/A�Ն�AV	�����2�H�s���
L �it��E�t�78g]8�_�;�ϯJ$ٿ����9����PT�Bj]�D��z٨e+;m[;��+�NX2g5Y�N�^H�t/N�a�F%��	Qi�SZ*����9ֲt��֛2+F����fWrB�-Q�����N��+g�C|B�V ����Z��*��Sӄ0qu�D.��f�;���vv��om�i��8x��+Sl�Ș�ߡ��{DT#�/���hsEͥ�cM�I��F�@�"Ka�ˇ�G��^�#���2t��Ԣ` ��G�8�a�Fw�9��ةwVPr�pJU��k�Z`����߽ ���/����MDHU �v�}Q��N����¹}�N�g�?${�v�s0}?�3A��$r"V�SZT���v���\��8���V-;ӆ@4aq��`1�^m%,�rO}�>E��F�F�a4K��7#�cu�Ro����%+�U'��|�~{�ϧ�5���ﳯ��u�Q��&D��q&z�L5��狇4P�����rUn�d���+.��s��nM�1mb������8\�%D#@.E�
�}*�F��n�jU�uQB@���'�t4��?�_��Z��k�f,T<�F��[��
Zbg���^�Q�`F����z�^����F��ai�܇��4Qz��<y�=����B�k}/�24�R�>�*:F�ǧ#��(��iJ<�����ұC'�P=g ���tάv�	()���qN݅�V-V�َ鍊R?�"��TlODӀ����Khm7Ld�+�~q#�p���>���ߣ��x�#�����.[�d��S���蜚�-}��9����!����n�_dE�����P_-o��d$���P�U�Y��{1�)E�v��'6�)\�
J&�:�.
�	�Ss�h�c	?��Vtu����R}^�8jm��]�6:ܘW���Jp=�U�`Xƫݓ�pXk�s�o��TC�+��D�-"X�N-$��+l��	��\�\�u̺uo��p[�G�Ֆ�B�����~ܸP��j9p�:Ĭ 9�*�C&�Ė�E����K���dTYY13�#yl�̫�
�I��LG��W��} Ð����6����w;�;�����e����s���=�a��HP���jS��0���H����#���f/n�n���>eh|+���ߏ�m����r]��,�pa��|���S�>����v�L2ˀ������c�l��ֳA8y"��A8�~l��ܖ��۸ę'H�/ �-}�����e��ыj�@Le��SM�	�b�4ٹXZ�=�~���g~!A\"!(�Td!Zl�b�'��-��ㆦ%���*!��_h���t0M�lQ�P]Hܶ�#s����UE1��_�M��k���9K�s�\̯�e	�K	֛�>�8��>Tp�����ǧ�B�,���%���%���=�5r�d���1;b�~���/i�ٱNn���J�h����t{ı���fI���'�y�v���pF�]=�$J2��'��>���T3�6���<��VR��>� ����C�UT�F�M+��8[��W�٘����U�69(�D����.@��^Ǡ���M�#�Z���lq(�&�y1����rz�)���I��IU�`���5�iը�ֶ�콚lowv7(P�}xx�Xz�'x��w�eo�;�t �m+�P�Gg�|�����r�ZP�rGa}���ǫ���G������Sb`>x�5yX��s8z�WԘ��gʋ)���/: �6ǋ�̃�W	NDwd��sZ�D��y���3�'�[�wK1?�bq��^��'$D�鴘#��
o6m�����E�Ra:1Z�$�S�s8�n�wKU�;����[�g��I*]�'*�:z3�RZ] ST���E��JO��l3暴��[�LRZ�M͎��^�./�-tͭM��@Ʌk�m��p��=~�����g�0��_Ǽ�v��3^g�؏a�Y ��Q����W�����78��@4�����jk�-S�)]o��G�=�
 N��PwZ<yWs�*�O%V���)�E��j���4j��YG����"{~�1�3�|+�^?*2����l�}"�^���LP{Q s\h�l3����߬���k�T�4s�j��`��q�9"�Dn,��:��Ǧ�"O_e��>"I�g�qS���&��8|��	�_���
�;
�?Jܒ'�u(f���M�$���9)t�t���H�.%�v^<��J'j���u5�~"E4/�����f$��7�p8�F���|�ݎ���˓��d�!BBw��I�.�ށ`��ؐf�H[�L��&��&�?��K���V�Yľ��6i�T�_�.z��Q�q�"�$�����=���*r�Gv� �t��Q���FP$4�x��}�?�%O�.I�#_��J�ř�b�I]ZM�;��3����?y�����)�#��_(�5�?y,p;m�� Ao���1��:VG���7�;'�+��H�����d5��x�+�D�ɞ���%���,Pu��e(�{66��@����~����e
�SX5��n%t循�m��4�u+�6{ZY�����Q0U�@�����o\��S]}⠧iz6�h�d���`�����N�Ɉ4����_F��"CL){&k�  .E���u��4��؆��eW���m�J��W���y�����Wiq�b-} |GG�A&	�Z(�V�)�O!&i(�r�U��
b�UnE�~,4jB1�?
�xg�@^��?���p0Ȗ�9U��K��zF��uh���M�9��ϓ��5�cV���G���(��Cۡ#���Y OMXM���ݴ7���nEs9�
�o�|ΰ��n��%�0<�xy1�F�-��GI2J"ቶD^�S�c7I�fc(gT�/ՙnY� ��RMw��a�JQ��e��`7o�%�VV|P��9V��u�)�_���
w�DOeF�FD�턅�Ef��v]D�� ��˭���.]Ilq09�c���b�����5g���N�e"'�|3w�`��4���L���� sj2u�3��K��~�8f�G%j��=G�����p�I �g��������!�?�io?�����j�a(�m�cVеB��_��d�uϋ�SÒ6!l(��g6R�E�ש�v���M_î7�)�I�Dk`G��?�]�Q�?���r�Q���\�E����9ކ���x<Jq��c��|$����!	��4�࿪�Vp�2Γ;������B��/�v��# i:��A"K�2��yk���Mz�\��6Ln�[a`���Ë�������ƞ,�8������
-`�"���厳dF����b1L�9u���������]9J��w(L ݜpe����M��(!bbЇ�Y���ע�4:�`rn�by"w�|"�;ש��<�b[X�V��rO/%����]<x�N�a�OS���W`g�ZgW'��a5k���iy����#�ߨ���2A+nE����6����~�N�X~3{A��ub��i_�M�����F�k�ݟ��gHJ�@�ZA���ċ�]���"iPƄT'���j���7�J���Į.0��b�h��J+k2�E����䟈B�?�z��U��S��د�l��oJs�L!�����m����V�Q�cE���@��^�E�E.�Ŀ6��!56����1(� f�^�̸b)�o�UQ�`8�{(CJ�ϸ~��ǟHs����6�
vU��c$�~q��NK��J���̙� m1���E��o�1R�6$qC�OH��-t��s�.G�`#�R���0�MӬ�|���}D�X(�
� ��B�#�m� h�@�g�6��	U�%�Iyy҆��&rW���ד�:	u�H�3�H�W��4C���vǴ�Uj~�?)]E��Uj$�ܬA's�B�ൊY�\�*�DC�FS��<�30���a~aGφ�6�U%����U�TY@�I�h)���*V�N�d�Y-�I�#)6R8���O���b��(v�=�?���^��~"I�g>�D۬J����T�Ʃ�Q��sb�D���"���x:��f%����cp˛J3�G¦�г�ˁo��|�L6g �`�,�����}���bRyn���T�=dnr�sF)d�fq1��|�U����s�'d	NŦ��Rh�4�=���x��P�eu�N$�����ͣ��pE�oU)�k�6k�1ꡜ�װ4�ãKw�-�,&�L*������c���LZ�i#�-o1�tq�؆�D�(C�G�[��X!�U7���|�iO0׊ԭoq��$�½��{4��s[��>B~�a��8Q(�:�p̦P��-�6��p���ҫ��Q.W`�j�/��cu$z,�g�!M��
e!U$�%�����6%��Ϙ��~��A���J�8��W��E'�IBIF�/�Z�%f�n$����^!����R=YS�C��������٥i� &a�pqe��}��s��dX�}��)�s�̇�1������j��Q*�13�8��z�@�vc���G���$&�S����8���\���	��d�]0��=+�[�S���-fy�5�h��Ƒn	T�<u�yH��u�U��!+�K
d�'2����-���p�ϭ�Sn�����l��Dr�~QF��V�e���W;٘�kb_6i�Uz�)9�0Px9�;Gix/�e��{��=s�5���ʤ����gñ�;v[4
˱}hh-]�g׮��U��t��:`W���M��pڅ\��9�#b�E	����{��`�@�|��'9f�3�>Gw��;ߑ��`������ ����SN���5�اK��|���7Y}�����;vQL	�n�f��W�}I�.��Ԡ0�6C�����c%�a�-C2���_N��Ba���q���(M"{1�d;�f�\Nڶj��+�i�e��
�SZ,
����[����f�e8�'&�ou�.;(b��;#A��H�����B�)�����p�Mb?��<q�ΣHԃ���8̫�"/��Qӵ�͘��B.�=����n�&��j�k}C� �d�^R�S��4m���"��yCSD��E�cX*8hz�?
^)�$��9y!:oh�S9��[a�gC�K3j;�����R.c��Y�V�,�L��r**v�r�2s��n�q=���O0V�ю*u|����ԝ=X���y�L����+�;l�#KJ�9�V��Ky��:�y���(\n��x�|���#k�:V]�r�5��Q�����vby�FبhvB-����`>Z)%��\�2�N���f���w��=̉N>����vΩ���|3r&�#��!�|�����ܷ��@�� ��l���q��<n3����Y7�.}�8�7���|�0L� �<��
��\ب�v�gr���������\CB|F�c�Y{�@���m���A�V�>�~	jV�Eك��jWg��Ъf^���<��=�y'g@��4�>x筚��V��h�{�A]ڈb��T+"t`��#zf�dL�4aY@���s/f<�Ks"�}��I�ڤ�by�&���$̰�^���Hv�h�a�y��׆eJ�7X��ʡ��f�A�>����%�H®�vyr��'R���q�e;b��\���'N�ݦ�(��)6pg������ǁ$�ލ5g��O����Bps1����#B�����,�RzZ��`����\Ӊ&0d�֯Fʍ$7cU+�p����_%R����:�0�����Je�ÐԶ����|�-��fz��lJ�|�м�ۋ-6R���w��r�����3j^ϞB�t�9!!M,��/3�	i��]���lL/f��z2汢F/�@�(��B���M�)6�|1fߠ���y�xV����P#b����#`- (��w�%�\1��t��\ ��Z��0�IC�nh�W�'�?T��!!�N�`B����-@�h7�˅�z���[ӓ��6���9��Ȱ���T�b+L4��:��:�j.�j�"��v<����6ho�Ǜ.�n���

qVɀ��;�2V���w���S�8�����Rr1f��_"G%� hyO�]��XC�C���@��GnR{yy� M@�{�
��ƮR�ܙ:�3d%/k�E>�w��1�^�Z9���{��*խUơ�o� +��ov�@�9���7�U�^F�n-������[��~��!?ν3�UoD��,�Zrj ��þSL��V����;&"ho��,����@@�'JF��q���"�L5��q�����-��mU�e��&ζ�G�}�C��t[+���l�N]Ɇ�nM�S`�b�u+�{�)�>٘�~Ɖ��Kd������=.m����xo��Ȝ.�|E�2 ��A��}O��H�PUv��qx�e�7�T����@}��/F�rAS�x����w��P@��l|�\f�jF�虴�6mN�	�-�6���6���,��L��+յ%g����>p��o�h:4����:k���Ȉ�ǣi9�$K��ߺ �%��]Oq4钒��d���'d�#�py�;�u4~A�-X�c��)��:#i�U��K$H8Eb^������Q��2'-��D)=���0��ؓX�қ(�.cH3	�p� Ǯ�@T������"�6�eє����V��jz��	���� A{��/<�5zgއ��QO�:��8<]��mk��f��� �w�c�F�C��&(�*rB����������č��x�),�]��}��|(�pg��j�;�'��y��1՜=7v�m�|��nu:<{tmF���^{�����[`�:���Ne��������B6[bs� d�9�W !��t%]D��Sb�Xߐ�I���S�c���2�h���������j.�Q4~�>�s1?���d��%��(^�S�4��|&�Z�P�w��m���I��5}Mb����Y)�����]�t���jW!w�r�*���T]ɋ9�O0��O�hَU����W�Ƣ}M��6�;���@�&Y�;���N�~2FS��hL-Z�UUi�%XQ����m.!��*�jL%��=h���Ӱ�b������k��E�lo��hl~`Tu�����(�}��xXwD"�P�0�e��!�����[?tPʡ#��Щ��e���ƣ�{V*�L��Cq�O,�8�4/���)�������b_�.��60	e���_%O�먿T���u��q��i���N�yy��\\�1Ā��7M�SvL�,D�i�)���={�Gl���}�|~�����An#��1�g:Aa�i����E�t���Y袇M�H�R��53_���h=@{o�s��azQ�>���\�#Pݛw�g��-��S�05&o$s�L^�.^Khk4�������7��ZX�� ���a�,1�=�2���[m���q�S��:���t-'B/ 
��ۣ��H_1Yo�z	ss����u��#~��d`�3D�]���8�.R�O-:�>[-����0q�gKO�Û<��d����� 3����%�(��u�j& ���:��ZO�,SU����p��~�n/�F�u#oP�S����)͈�L��ݿ�e�H4Udqh܀(�7O���}�*.NDF�^�.����5������W����p�	J#��2�l�¦�s(4͟���0�8 rF�\������AZ5O�^��K|����L�6~�^�%�f�;����$M-Da#ď�|;��~`����k��nބ?4�[� ��3N����U��������[-��
0@�Q�j�P�B���= os��O��q�9\�?lvڂ�㛚��6��i��ܟ�^�=}V���3��oKޱ��,V���{B����a��?�ZgjR�b���9��w�8w2�,��"�/>������nn�}|	�"Yqh�5���8��x�dP��y�$����FP�Y�"�n��ťѬKv��I�\�(�FoA�dJ�%\�$��ۇ�[8~��|>;~��J��6@�`^R�q�X�}���܁�z����j�iS����g��;�"8����T�hyȼI����G�$h '�/����`M	
�Pj;-wYqw�4��~���"����d�v�Y������s8��Z��^tc��`�6���/m6��V��'��`1����=a
�4�DY��\3��x��-��I�g̽�+,N�?��VÿP�B�@���;��q3��a3OQ����e���B��N�p7���I���!@s���YB=���л�ƈG�D��7o��<�-7��#I+?�gj�2����i"�Ok�Ou�x��0ܖ���kvA�ϾCN~ʟ5W�bf�����O����pZ~^m'���=%���>���hn(NW9�������(�,��ܕ�!�m�>�Y�_���{�'�H9��D875/bD�ŶǑ�l��!,X��aHR@�)'x��B��B�IQ�xNg[TT*o�me65ԝ����dd�������fF�qP�U�=����ă角E&��`^�v��=��=�9~(C��E�}��+�{D8��m�4����rUrU��c���*h�b��["׭y�j��3$Ĭ�(a�_Zg�G�s��� ��Ú�G	�h�^�'+d�d�q-��P��A��&6����P���=R3�o�]��3����z@ga�֌A��҃�1U�~f!�,�I�@\+���-w@9r�!*|�����T@���!��9�S}2���Y�;UA�Cjh`v�ږ7�h6�k%�T���Ԋ��d~�� C�ekؖ�a�� �H�6Ώ'3{��L��U��t��Ɠ~�|�t�r,'Si6�SW�D$�U�2czmc��}��4������^�(�A������a�R��CƷ�g�\�o'
�%u��j�z�>��Y�Sh9/�T,i���{2�	� �J�A��!w�x�ɕ
 ���A��/�\Y���úy��¯s<�^�b��l1U�y�����N�"����NҤ9�&r2yF�Yĥ+�:��uO��"v�J�����m�w�ny	؝6�W�d�yT�w�>ۑ'e�j�QCL�U>#L=q%�z��*Ei�%�d��2��af()U���\_.G�6�����vBz$�H��_�2��Ϻd���?��XQ�G�Xm\M7)���\D���Xz����y��)Rb.|d�]ul��i�z� ��_<��.!L��K?7[���C�����Ono� �eH��4�>�ճ������o������|�͓���w���0��>ao Z4ə��ृ3�̓����oN��X�>�SnK3JPq_�i��u�w=�N��ˬ�6f�AE���x�LW��(�O��(T�}]���������E8�f�m����f��ا��E"d�w���� �-p�}4���A�3g�[�!��~X˺L��Gͫ3a������, ���?u�`�S����B�~9re���7f�!�
�K�P������:�5�of~�[�
���d �2a��p;,��%v��%���]5P�� �T����w�GǣPg�>�Y��R���13M����SӾ�'R����J��Ym��/��� `���2$]��ɉ��L�.��:v�h�PM���^;�P���&�d�����|]�*�'�Ű�Y�m/�ʩ�"2��ǿ&�!��~��j�	XMе$)�+y��m=�5�Ԃ
U�6��ʚ�*	�'R-rL�O��Ss��C/�y)�8H��*�@�┖��>��y�&h'j��L��	N���)B�{�0ǂ��66V��q�?̞ q~QG�SiD#XN�Ǜ&�/hh8W�&�Xi_!C�ㄖpy�nϼf� `�_$���N��y}
Щ�����:��a���O.x����9���L>6�ˁz�x�}�C��J���
^��#	��ۜ �9�$�=���q��-�1�����L��rD]���T�P��$F�fd� �)��ڟ�n�:�5�����8��=�X�r⻖yg�bs�Y�qY�H�qJ$S<��������7���@��}2�>�Q����3�!�� ���J�S��?Gᖭc��w"G�*���&�b�T�@�R�"*�t�Ӡ���FW&S}.]�]�1��c*����R�YQQ8ah�V��Q�+)�5�s�vl�:�"�R-�礙ټޣ�L_��gO##8?҈��#�ZQ�|Z�ϤX�[,~����cm�8+Uq�Y�I{C2E�zv����`e�>O��Ю����:�&k.8��� ��%�+�o�[&�e"=&�.p��X�*L���&	bz	U1��m_I���Zd�e�Xj�+֝Unݘ9�	a�����DXw�H�(�j����Į}���塡���aM�qnJzC��y�?^(��׿0���H`�ؑe�j�-S[�����Y�5���������!��s����k�X"��˛����	,�U/s�K�[��u6(ͣ0Фk1,}�}�0�Z�6 ��H��Ɠ��@Z�и�
Y�
tYk��؟�^�4s���&�����\7\�B� 0�Y���"> z�- �5q����+��:ۢ,�T�LH�.��&@nyl����	<d�9ݚ�{Q����Q=�lɱ�;V[�HM{r��V�����f*�]8�/ϣ�W�?x���{P��fâ�Gi�����J�̜W�z�p�a�:����	�����
Sg�� Z,�;�}^�ڕ���=�T���N{N����'�Ha�7�g�f�S�wN@��fK7�i:l)���������������p�7���w��i?_O�+R�f���{�@���rGMO7��vL�{��"g>��z(�Lo��(9��5#fg��-Fbr�%J���vFg��=��Z�UY��U�?�����*��*p�oW>*ZH��DX��^���N�y�$n1��m��:��ӫLAYFB�rȮb��yk�����J�����չ��f�b����~V~���{��ML�ze��d�Q��\�&p�};��(���Z�]��z�����S����� ���4	�X�i�������ϯ(�Iټ=������S?PBu��^Ф����$��P�>�ŅZG*H�U(�R���͛
k����2}Y��-G9z��e&��61���
&�F��r��|�����xQ�w��	���B[�����Ck���">)IcR����~�����^��QNj�C���Ӕ�q�Ӌk7}'h!��+/��1@שק/���cFw��P��x�'�
L���`+��&����e��|>rd�Fcܵ,��Ǧ��1f�aI�u�I�4jD�ϛu{�Ex���� ����צį�yJ��Z�o�0h�}�3�R0E���X���z침��<Ց�1����B�+v���1��H��E�C���_�`��u�����o��q��X�~��� ٵ��p��L
���S^%sk�i�:���#�J�~t���,��� �*CeYB�� ��i!��u�9
>�U-UI��n��'��Ɣm��CK��d���� �&��xJp�����9�]�VZ�o�2���tUq'����K����=d�?s�T���z8�i�d��4�kz�\�zx��<���5�rpBgB�n�2��M	�0TY�m���XS�9VrV~Dᚷ[kJS�8�l��<_�^��9��7?��m�A�/�Ī�RQj<i���ދ#ՠv��ӓ'�Ѣ�BH���b����΃����'3x'R�(Wj�b$H� 8G�(*_<7doq�%v�;%�� �c��g�4���m��B�o�o��佯��v���L���D�.�F�3%�DSI�	@F�����2�^'�O>Fsό'|��1��F��l�)�m�.�+�!Lk��9%t��;G�؁��I����]���j�{��F\٦%>̘��-v휛���~	���Q*��c�0Y�"�`'�,���A���i~FĶ�0E ����S��#��1�o�t�x��=5�/�Q��Q��� �`�yP��GȲ}�l�ܩe�K��X�=�O���v<�j��B�&}hC5νe��i�Di��a�g�f 
�n�����=�yψSB����?[Z�[�\S�;þĔ�����ksѡ6+2= ���q��N��OHچ��yV<�֯[Al�B�y  �����'�y�bܠqÖR������⮣�����[*]�8͛K�l���Ka�>_��Z��@��g7�`^1����]I�1��P��Cȓ��[��k��l�Io"��i�;��w(������C%�ٛ	⿓:�������~�6��f��ϤMi
Z�Fb[]Zˎũ� ��%W��"��/�\��=F�M��Nt��%����H���҉�=GH�V�4��x_��hm�Pk����j�	��$ܰ��&Z�<O���~��r�v�r<����`.Qy��3�`�J0�[���W�Y�ތ�
��`e,���P����>��q���R�ku�)��|߰G�j�
�Xtb�Gz>��ì�!>�r.�wx,_k
3
R���C@��IZx�����^���b�(�3L��Ͼ4A@ ^]���|(S���rtå��5���B�ކbB���6��_��Dl����;�����~~��\��7�)Ni�Ә���U?r�'�>C���
[W�+Q��4l}��BL��E����M=�Y+�A�s?Bf/M�nge[X�l�b{�lպ!
]�.�e���؂஭B�ہ;��-_4rx7ɼRj"��͔����쌼zl]�@�	:��ʼw8��}ڧ���{�t*e�Dq3��%��T2��0g��n�
q����ιy� `-lCȕ4��I������c�/���֫c$BV3�@J����k��d>ǥ���I��d4n��N��;֋D��;���GO%YPD��9�"���-���߆�K'NM@�`$1ސ��eDʬ p男>p��h����L1i�����Bj�1S�L� �0Y�P��j[�
����\�R�L�~j��I�$x"��y��l��o�PE��S[ ��=	�=a�e#i�I�\*�߮���}�%`1́�>O�%�E�l�Hi��,���(���=l ��S�ޣ��X{N����y��N�KK��w�~�:�tcL����H��-�is����O�mZ<J+�#G11�k$-G�AN����玀J���u�?�4�����z��`D �(a��g:�z��7[$��.V����D�ѯ���R=����cו5'i�T���cA�lq>UI�/�*��T�j�m����v���dS���TS�?��s;����~x��X�$b��@�Q��$8�����τR��MƟ �0���9��h5	�>�\2�V�<��Snੑ��;��M�wR�%B8�S}�=ῦ쉮��������1�o���ˆ��ԝ�Ũn�[н���t�h7�6Ő"������_�V����NEb)O��S����t���^^���tdN<Id���y�*��Q*�>���z2�ڐl#`��lbHҎ���Cc8�Ц0���'VHˑ���V� �,hrD�%J�m`��;�aC��tJ��*�q桗�6��r"��"Tf�H$�{���+<�.+�gQe&�.��֒�/y�Yp?Wm��6k/���Y�َ�<L��Ùc��Ǚ.��ݜأ\cyn�����4oª���0���oW��Jx��K���c��;0�1�d���ґL��
֭�u��*�X�HX�Z��f�=�W|M
r�'�^��̀;��w���?e&�3{8�`Q�&0`|��>{R�����9ܘR���8e����n�Z�<����s{��:պ���cw`�lgb�Z��3�#qv���uzEO[a�׈���a I?A?B�TzG�*P�hw�{������#��_�I��N������%��c���r(��
;W��)$�i��Ӑ�z;�d��*�����'�Rjj2���]��f[�N�J�&�#��H���'��ǡ��X���?�N0p1un?	��2�9�ƎN�΁���hT�����i�e?_ E��}� BG�e#V�$%^��z#[y�	aV�Є~����GJK������]�F��t���2����B�1fK.�2�N�r������?M��M��B�l'�6Ic�1.7'z#��퍞�x�gEK�8,=�E6|���?f!`�Z�l ���\-	�_�f�*�e��fo������M�E�Lhi���P[��d�q�0?�R#*�S��#�ڒ��g�xT��OaH���ť_T=��E���Ilb� �utԝ���_����*�߰(-?P�0��U�������tTM��|Q|#�,ͦ��}X���������q}���f{p�b�*��ut�N��W����xJGpB˪�����R&�h��w�W�d�S�z��8�|ӚPhza�~�f"9y�{(u<@KF/�J
���4���5̩n<n	� �'i��K�mɦ^n�·�9R	�^�Z*)��Z�5؉s\�8�=�? ,|�o��s�yf���,z�ay�wU�Ӆ�o��H�蔂�2~��e_<đ
�P��7�Abvl���R�b���������l7�AW�L��(�������-(��fA'HD����{r}�'n)�D.�ļ2�-�'�(����Gms+���!���=�7U�[�_��=�cd�H1v�?�罡όHL�'��F6�	�����Lj)�A9�(�ɧ!l9��0���T��Wm���������i��uᳺ�/Z����k��Q�T��P�I*�� L&�� 渽h鲉R/T/ H���&5����D]>$9@Ùt�yWc8=�@�`V�jf�,��Ōt��$R�o ���	ܘY�����R��s�N/�W�����Co�Θ�7�ٸ4�j	�UW5�6��J 6g�͍����@�Jql߃'���_�j��j��N^s�{j������n�U�S����`�Ou�1�ڑ��v����/��kAV�WzpJ�ϥ���N��k4ɸ2ۺ�O-��y�P��y�� Bڮb}J�X~�I|�Βe �˒=�O��	�q����܅���;F&$���v#D(�\�2����e�VND6����ه������%in�|������K���s��;���xt��fl��M3tcB+峩|*��"&���#�Ƀ#��^ŏ���{�ְ|�0�5��z��܌��m����C"�wZ&��k�}�Ej���ż�'0���A��wX��A'��D��R3�*�ע�Eڴ�%2e0�%��[~-�t  �4�4j�f���c�]9�HS�%�ħY�B>�|�(wԔ��hܑ�4T�l�a��|9;��U�����C�	�;����HZ�@���	ng9h^a�,�j7�WF���|��?�E��8#M&�R��2x�>at�!����3�:)e��SSZQGD�`�sk�,/�yC�PHB�GgV�� �o�#ܚ^!�0?:J�|
��`�	����:Elw|r���`�+y����]���LŮ�*Af�;{<cg	��q��i����lU���qЌ�|���R���1����ןCWS����-!�LZp�����ʖ���Zu1g�qH��?kڧ��YFCɌ֟e��q~�J�9��|��o�éB���C3��x7���|dXX.�yv:";�
�ԋ)4=l�w��c�S}�S�v7�٘�o*0�v_�fD�
<�]���Y$�����i��i^��,���r&e tJ��!zݫ���9S�㛻��CP�n���}p�k��V@K1�����ӵ��a��5�Kȶ�k ]�b"��[o?e�vf��5����,�Οl@R�<~`y��&���^]��� 8�jN��ݻps��ү]"��yD��D�*~CA�na'n٘w��D\<����@8}Ow7��;6o��KD�����<<�����9 P9+�ZZ�/�hO���͵k�����!o�$�Q_ƣ��� ��ڳ�P�^��IaIh�G_��E��m� j�s�:~�ʡ��l/�@4)��U�����^��膵\Pū
��m��5D�%\�i���=7����AG�(J����Tz�,V,��\��#7�(�6�����M���s
�ݗ�[���/-���U�$��FL��.f�R4�+Uq1�M���5q��ME�� Hc4}���[\@k��f���P����Q�M��W56j�7�&R����BK-μ��uEC�E��A�ҧS�q��%'�"��	3~���'=���0��
�3M[SU�Î��RC�gN�zdaX����o@�8�#z�ڪ����i��J����K}��y�gO�5f8x'ҝ�����5�N�EFݮ+j�!	�K�4��O��%���w��:�P��A����&�?JZ�SӋk��1攝A����9�n"@���$����WˑP��]<�P�L�����`��$�s���R��6|d��p������oK�v+����2N���nY^��o�ʳK���}Kb��^Le�Qk�9��f��\��l3+mIϴ����o�Ĭe=Z��m�}�?��7&��h���`�O�d����@��x��o�+m�gl+&�'�9�a�bd4Q�ۈ�e�g�����Ż֕R��̰\&��o/���$p>�_Ͳ
�_�T�?�}�ަfu�s�-�b�C-%����'$.�S�t�AO|�@�<Z�9���[���"-Z	���8�F�W���k����X_����� ��spq����� i+�Fk�	����1JB�:<WJ(�k�����0#.�ǰI�p�,��\u)ڨY7�U���b��ph��IČ5��O��	�l5�|my}3b�OT@_5H�#��-��l�;;]��;~��\>9��}cy%J����5a����ڊ(�_q8~gd6��#� ��Rŕ��E3��	�P��p�8�#��UUd��~nN.��bv���H/+��yt��� ��ő���N��<E/ȫ�8S)7�bZ��o��*�!6�Ɩ�'ф����V�Qv�����K	$�tƺ����� �&F#�k�ܛ�j���'ݔS�K���%�=Į��n�IO�tl��s-I�|�`s>�)0���7���R!��Ȋt���]$+kt	t��
 -ܻ�rg�L��k��KqX�t�Y2;�B�5wk�~6��-��� ,d ��-GN$Ў�����	B>����#��*g�H`L���-afK�k������Y���M��C[�T_��Ȃ����w`�W�h��c�p�IL!�˯]��$$֗��˫��3I�t�����o6vc�$���Ŝ;$�X��L�\2�89H�Ϥ �,��>���(�c��u�\�`��������SG�[ ����4'�o�/��r���+��?����^죍�i]�/F.%���WB&�bd?F�O��d���H�����~�@�A��|�&��z�9����֥�N[�[V����#��������1���Yd����8zGc�I�#b���}\O�X
�]���h�7D6SV���Tc�i�}Ɲz���&x7���죌��N��a�mQ����)���h;C���������踆�!������'��4�E�L$ԡd@�/��I��7��I��ׅ�=��N�k�����ĺa��N�Pf\��ݳ.+P���ǭ�LDN�s��W�6��n�F�{@�w������L���#V���I{[#);�UI^�)���H)�Q�g������$F��w�;��t�ԧ9�%�^ Y�����Ò-QF�
��=t���%�*���n����G��&w��U�~�`��E�uW�c�xb܄�n�H��A�A�M�GY��8�Ϫ �
�#�zD���z�)Hw}�R�#ҵ�a�}�{@�'B1�g�[Σ|c�E&쪑§�G7 �?q�ty�� ��N�x�}ʚ�d	n�CYbQ8�j�D�0���9o����HE�P 7̨�wB��&&_d1��DK�읠̇������7�:��Kl�w�'��xMV//�$"aڻ���'�!
�#�����v����U*���-���2�n�u;��/[g�0�]C�8.�q��X�S05W������d5XAv�-�h��W���9�fJz�(�8�s氱o/PG؃fߒ�!h�1��Š�9������@?��tL���~@mņ���͸�Ul���(�04������!�����4��G+��A��IFRk���d(�>�&h���)�?�g1l���Q� `Sh)�,b����dT�9�xt\�j�h:���P�'UM	*ͫ�`��Y�4���]��ڗg2ʌ�����Ћ���ӓ�x ~�[�]�0{�K����R!���@�K��}�o �Ͷ��4G��@��Ut�E��"]�1S
	P�jM��7�,��-n����=Ƙ����C=O���P���.#Ζ�ծ�G�!"���*b�<��)�ܾ@�E���e|Sn"S=�Ȗ��E9;m^r�}3�s7��*�⒯���{���s�?͒	JZE�7_�hґL#P^:o�ձ����O�L�:�N��f�^�sv5��f����E���� Sd�"0��Ou�p={��L��0�߂;fc>�q�Uw��P��e�o��۶֪k�,��y7;.(�o�us���,���c�uŖW�#,K����ڕ"�An[�rNۚ��TM\��.k�h����WL58�!W�C�W���a1�~J	9�Y�=-�j��Fr"����ka�<�ҵ�\9,slF���
�.�s9�4��i|�&���6-�{͌D��V�d��D�R��!���J�I��[���ceqsY��:82Տ��,�$�9ubvf��TZ�~L�^��dӥD�n3� �}Y���Q.�Ӕ����L.�[�A��%̧�dTZOۊ��O�����0�3FS~�]��12�҈���I���0L��ť���l�{c� '�iBs�д)��~�v��o�h��\���u����Cy���H�R�^1y�Hd	Ґ��\��)���!�_����i9O6�&a4:y���c�?�f�Zl<w��9$̠B����hQ9K���S3w���v�s�R�4�;��ّ��Z�9�R�Î<�e�"���2����ሴoYL��N	��,�" p` ��"Q,`�q�
���O�-���Sy�Y��<����<Ĺ$W�7����(c���}jZq�_NM�]�#����-%25���"�z�u��+w�#i�RzL�kJ�fu���b����td�%o��qj/?�b]��+oy�H����/P�������0)Ȭ�z(QM�:�	w������4#|V��['�r�����:~GxS���c�X\
����b�$��X�?�R�v��Ù�9��B��^5�E�ՠ��� d7�
O��Y�h�AF.'\���W���]�@"���Te���?���y�,2�LB5�Թ�	�-]-ҋ��td�ٜ��Ϸ����>"�h�Xj ��"�bq�$.�h�"�%Q2qX�G&W �<wb��W��b<V5�SGΎm��H��|.�R�*r��ǜ��3��6̿����o,�HC��C�遺R�vJ�p`�
2���$���b`(?��������ď�v�V}�[��\�z�g'D*î��n[�3�~�D���<�����e��i�u�P�;���
k�ʥw�0�����y����;m*E�bM�����\�2+���^j��W Oƕ8G�)H�~a�q1��!��	��7���,�4R�eh�Ii Q��#�M�%�W+�3�_?U���.�`V�f��VF������;ڗ4��t�[�+�^�f��e4Z���}l+�a�%7��R/EtVw�������F��:��$��LX�������+�թ��I��T��4"���:Zԍ���o/��;��ݷ+^1����;	�-�759��Sѵ���7+�)C��*s\���+��u�e��l:_M�s�aŉ;��3���lY�ߡN܏*�ܐ��sn>��ĝdV�)k|-�)?�-"K�mB�OD5o8X��� ��А�r��&^%�a)�6�-i7����9C+B������o���|ͫ.Ü=����9��Qz� c���ԫ��J8{W� �Y{�C�kY�� �
��>~C��@Ƭff�K<��n�K1~�ac�(��������w��k۔d���j�ְ���<R�Y�8��F��Y=�qɯ��X)�#( ��r��TIT� fpR@�#7N��㬅,a��86��V�������Ob�J�Z�({�7�{q���W1��d48ܞ�jeV�P���r���tS�dg�n	T���ӏ�tɒHi���Bm��ms��P�i^ u�m�����<d�B!�X݃K���(��߲�U��ĝ��(�D��=�]tmb>�i�8�"�7TVf��H��3�~�@����;oL�o�"�B�ē¡�W�P�N��`�A\)�Ƣ�r�[a�[�e�'���|��ʨCv����9-0	ᚑ`V����(DrD\ţ�<A���tg�zG�T�3���?$��9���:p$����|B�-k�ԗ�T���K}�
�6��X[ԅ�X�#{@�g�|��DK�Sy&��@������`*�Bf]�� ڒ0pv^6���w,���m���3���s�l�񦽫�ӻV�p=�`�鼑���k}ف/6�8O�Q�Ц%?4:�����[N����_M���av�t�����V�;��Z/��k-���d�[�p��ҝ5�����T������t�����t�8asc�4��6u�.|tb��t[�B��w m6q��������VN�47���wqIΙ�wn@����=��ڋ�B0ËaTT�"��MM�e�A
��l��B�`��,��xfYۨ��Yn7����T���u���5��=1R��4r�i�ɋ7���� ;�h9	n�5ao|/(��^nb.q�_g������pe�-���ו�_����� k�s�.��Xʴ��)�*u�Xj�>�Ss��CU��;�%=k�
'�n�it�d+�����M�͐��+�50ր���e� ΂����)9�de�T�+��=����?����6�X[���MZ��@��f����@<�Vr=e
.�ث	��WÏ�x����M�d0D�h�:t�8�&�֭N�T��Y�*Q{��n��]4��;� 6wĸ���B�6�?�w/Q�8���#�o/�ʒ��G���"�/}<�?(�F��Y!��}���Q.�@c+G,������)nJ<���W�ݟ���͘�A�;��+���P�F����x�������R:f����Hݚ?^�&��0w�*�����hU�-㺙���ixz̆�@儜ĸՈ�}��~����B#0B�6�����)�AX�(��-=�{���(���;_h_v��D{���5[�Y�vSTn��v�z���1�>�SF>��(A�3uVS-^iP'2��Ӿb;��>X.F�
)(���6�u���H���u�+�� �*5�:>yо鋐v+��s����6�w��a"�͓j5��1B������J�k�]=��x�
9p�V�8Y��QtG8|϶�c���͙n�`�w� ݄��>H�����ѵ{CW299_�&���;�&��1 �v���q���^-����?	��(h�J#ry����p�K�醖�}��κ�����X�X��/n��9R֭73B*��(��`B���5� �o*{�߃{f���bY��X���>H�m 
�`�	V���~�Z<���$�M�ܙ���(�|h�~��������fǯ�������C��̚#�<��>�b��]zm���L;��oe�����3�B�՟S�j�U���z�Pd�%o�4���e���$\V��\�V���$���F�|�E�N/է¹�<Ĩ_���F��l�x��9�WY�U��Sh]N�E��z�c�LI{���={"���/�G�X:h9C�\ŋٟ���Mf��<;�wϟ����4�5�i�X���
rY�.���R�v}�3ߎ����ې�8&�{�
{ן�]� *�V�="���3(u�A;�$�]�dw���ċ�I�@�m��(\�	�o*�$j~و��5R��Ņ���k1����K\���sX����U(���֯�*��͛>��< ����@��q%2s�2�]48H`�3�l��Na��)��a��^�z�b����\fb�b�Ӎ��=�Bq2k2y�����\�R�
�{�I��R8�ǖ�.% �/��v
��T>���aKu�ۗ�Q�e���Ǻ����ٯ״ӗ�����Bʡ�Q��$�u6`�������g��z���Ƣ�72hc,�����U������`�ovu������'��k��7g$��mv~�����]~�ʭ���P�G�jF�FK���3<h����"�t�0��(Lp�����+_2�y!�ChH=ڐF�Z.{��<��8D� |ˀ���������dh�XJ�=��zv��f,r�#�cgac�VP�D�d� �p�!�"��R5f�I<�(���=y��lq�]Ir������lQ�p�\AؑT-�.��Čʯ��j9���h��h|��}����g��z �]�L�Ϫ��P)�������������3����-kq�TU1PS-Hd�� r� �]?T�vI�s�Ƹ�@ ��s�@_xk_��Ϟ�G�T�i�V @Q}�RC���\o5�G�[3�)�����,^�C����'`�o�4Ƞ�1N���Լl�$�֤�����9��sW�qk�PH���T�:�o��Z&�wbjH~��;��>�$|�
�I'��8"Xh����)nx{=c�~��/X��n1��J�\&>2\%*	sd>�ה�J��b�����-8X� �u����Z?����7R5|�@Ӥ[��zj��+:Ԏ�S�>��[ԫ"�B0��q�uG��)��9��n�C����X� 
��h��) 0T�[BdB6C��/}���ˢ+6��/f��$
�|`�e�,��q�P|���R��T����F�T'��j�����fT���f5�#X����-	T
mt8�Ffu2vwpg�W�yd��c�9Y2�:j��SJ�A2�I�K������h�;{ڐg���f�f�૵C[�N�a�F���۝���٭M�0�Z�xqi�� }'�H��ꮐ���F=�Q�f�nhc�ˆS���w�xOJ@�X����<*�G��*Lh����a^V>_Fx߬%
2�s��� ݤ��KH}��	���F��@�P����ޒ�	]�5ܮ�˯��R/!~/���S��@
�g�F���D�T�u�� pN玂9��#bg��֭z����=p�"4X`��P!I���!����hD�Lu�R�j�c�6��J0�����>�O�%�*E�0������#.���H��":�G����A���@�����z��!.e�#Z�H�%�����@J��4 :������۵��ߒ����V�8�O��X���v1m�:�	��q���	MD�t ���?�J��)�ݑ���2�����4Vip�*�0�e�T��9��^H�="4�1��j|����lZ�Fn��b���������@��K��:X"�0��F�պEB� G���B��ɘ��-[���/��P��d�sЁ�\�]��U��e��Y=���(͜��#0�jlt�1��_�虏6�q3j�X�(xO`���;{hn�u��e��$�	t��x�_�k���"Lǵ[�a��o�C���[�.J��P���R����n�Hx�9�>D9�ῇ�F�q<�2�eFW���*��n���3��VQGûT�y+U98��-��W�e��֋�}�ـYK�������
�x�_VÍeqf_�׈Ӻ���ٛڨO9����;!�<&Y������������H��3��T��H���xƤh��ڵe��C��a��ژ.�;h��f�ف��}���w�Drh�R]Ԇ�bc�[��%�Y^r���P�;WQ��O�����@{l�8�Q�×��;| ��p�g���b8Q�v��BkS2|y$4����m�]\Dt2�ꁝ��Hjv�~���Aw���.��dV��r̹)kֺ���:���t?�2�4 ޜ�_��.�Q�wJ�rB7�
�7}4����2lH�P2�5�m���G���+;��@�+�ū�8���li��&K�̤�V<�T��Ri�s��,��#�A+ã��`7]��P�9�]��D�qb�oupsa��a�͠�2��>ϊ��<�i5a�Yb�������	��Ω��"E�����)�����n�v����ގ�693�M[EMt��/A�~#M����B	�QRZp�'Kv����u���PFݨщ�;^��GFh�qU/����A�
K.2-h>;8��;Mk��tq�<l����	v,v�F��������~"�nl���>������ԯwu����#H�q�,�w�0!�X�u�L���`��.Ql��^z¶T��0�,����H-Y6�#�!�kz��+p`2]�"�;G���\w�ŵY����b�N�\�Gr��$��6ѱ�����,J )3�i>�z,u��wkBw
t�8�c6��w3�H�=�P(���KĻ�@����|i����H��A9�z8޶T�/��^��ʨ�OʙDƪ����V�� ��MHP}���])��LC�S��
���n�e>4u���)^�:=ԖD�X��!�-�#���v��&;;��ɼX:����`�.U?��tƵ�	�o�H)�S�m����x}�K�#ܡ,ue�N�T�/�L����͈��0 �Hc5ܝ�����KD�jܡ����X� 8��&���Hq�¹�s� R�{��C0h�8`�w���s� �s���7��3oT3x����;�NR���Qv����F��&Z�U�˦!�`��4��\�v[;�w�/]2����q�=�C�J�R��K������A��q���Ҕ�Mu�v��O���i�*�s�ls_O��w���Z�mf�B�M8�F���M��J���vݪ����(=2�����' ����p^WdR���ᄳ�� ߲���R�Ī�q>R� M��o�+޳a��.��E����ΥM;��J��&�v>e��jdz^Iuqm}��{q��ӛ�\bE����qۀ���,^�P�k6Gꇴ�a)�E��ðݨ��Ө��+�k��*��XvԌxu�Q�ca���=H�����8P(��hv��Z�ĵ"�����\�Ϫ�H��Ș�	q��g[R��Ȑ��!��C�p�ϓ�qP�z(P��	�Z���Q{�)�j������4u����]�s�/!�! FS��Y��V�6�V\�O��طy�_�'��q��3H"=�t&��J�����A�]#�ks��iE�q���f�J]����>r�"E�2XYA���>�������|ӗĀ�Z�3�eK{�*$�+xu\X��d�Qr#����κۋ6b
�
B���s;���I���V[�5��Ϯ�g{k!ذw��{0�k/�� ���4��Ê�m}���$��(����3��(Q���%k ��_%_#DG��c'yߧ�2�]�}�0]'Wd6ǯ󝞲�&b����X[G��/g���E ����M�߯c��?5�3_|��Ykdp�XW-1d#�ձ�V�WzES�ˑ����h��L *��:�c�9�m���qKłO�d�X��[�"r����,%����e J�yY��'Dv^S&�	è�ݧܮJ)���Ծ�x���P-y��,fWzщ�gm�?�wK�}QU>��ф>���,|�M�@Mufj�\G�����_$��z�Q�'qx��1�T��\a�1n����߅r�%>7�`[��zFK:�e�<��	�c��I��gn=@��A��!������ޱ��Pt,h�v�6���(R���y������m��1���j���.��[�7 �\ ϕ�/	�u��v����"_f���/�.2���ۚ��RjVJ�w�2���9�@<�Q��1d�f\���ظQ<{��/e���c~.U�fX���|&�P�0�zM�A H��5���������2yE�r��*��^L>.�znx{{��2�9Nx y��ۉ��ǽ����$G�j�9P0�E��S����x('a����,��1��Ѧ.w\��Ix�P̨�2Z8}>j�X�q��9ԍ�g�cG3�����x8�CI��S�U��5�u N.���=L�$�G�U2}��N�Vq}�j�C�V�X�N���wC�]�
ل�,c!u?U��ڪ���I�lxD3/`
���[�W�:�����jjL�|�+���	i���a�#�,#rcHL��h])C��E�D(�����*Ω�� |3�(AY8�V=-W���Rl�\�y�ڪ���N�nCD��:�v�o�5�-��}w����w��[�]�9�_����H�ZZ��Ǥ:.�D�=�%~h�?���~�:�nN�i ��n���*YQ�ם�BMu�Q2S�T�l(�㎂�nY���"Sz�.M�x���#�
7��/�z�%���Řؗ�|q>M��k��_�r �#��S`x���)�����s��G�����)QHm���El���*��bO�ႛw+���9��v��)� j;[1��P�,_,a������LS�����iH�I��j+-�^�'�MkRi���1�f�4�LR[ .!�%�h��l�ϋ�Q��`N�?C�5���@%Zi�w�Zڭ!ՙ�VHׅs�"�]q�fۃ-�ȯ˰uQ��	7�&=�y'<�s�X��呝%��t� 8@�b��6�4�$S��v��6� �������)~S\��/�l�S1O\a���z#=S+���@cR������h�}���Le�#}�!�p^��� >.u�	F�Ҙ��^fSy�\*PO���:EOS�	`q>��A�)�0�0�k���b߃E\��S_����d��X���x+�ȰY���˫����Eh1�_(�^���7Za�A������ܯ歾�Q���&4#�8�E �"C?lK�;�E��]�60��Bq�� z�1QJ�X�E`��@�����Y�#/���5��fb���|��s�܋��|α��7j��T��_Ҡ�n<�]7�,�vR�c���*�xw�h^b}b�t��Yo6�9Eo"O����#3<���Y��ci�	(ݑ����H;xTS�lTXk�ĭa )��3fW�p��V����S��$ų7E|���[�ͅ��9�2}�bD�Zp�V�>���-~S�,a�v��r�LA�v3$�w�CR��s�Gtr%��u�,�G�H�u��M�]Ox
���Ã�k�TD"	�F��i���q�q�Ν������~ɅJ;B*�Ւ��o�Z�;˶�Zq�nF�l�D��-���Β1g��@.�~���
�M�jI3�ru|@�[<7��,�.��Գ*o^nG~Hf��1��HPy~�ӛ�
��q�Y�P�ʘ���*���'P��l `"��QK�<��*ؾ������[_��������p�9�:ey������+E,��5_��+����X�I��+j.�#��v赵y݌�e��3Q�-݀�ZX��R9L7͉��oU��e�m�O]�z��l��0�bI�3I{��Є���v��n�;���q�.��{�h��M)S�Ъ� J���ܛ��1���i���_(��#��� 49ǜ������X��E~q`J�k��c�+9ù�h��̕��߶DZ��we��(�E���aJ�}�0_�P��R��������s�M�Gg-�*�6!o�O\럊T`I��K�;��?���V�l���Q��e$�FQ�@H����oi��2K�!��EYE���ۺ&#�'���O�1i��L#���&~L6��H��U@����[��_�ڡ���GF�v�k��(��k	�$�+|nn�buQ(3�&�!�}��,?X&�����+(���כֿ�"K��*�-!DM���	I�ݖ��� �,���p:V��v�6
��
š#$�O�+��SK"ma�!ߚ�W�M�]SZ�	X�$W卼��t�k WY��X�o�a����Nb�~�o�߃e�%f�$�*�+�~4�X��n��c�ږ��WA�ay�6�����K�έ�g+6'�V0dߺ֧W����>�Է�t3��Q�ۑ��r4u�ݿ��UX��n6�&�
���O߳䪂)2��b�^��6p�L���z�F.�J�#�/yq�������?���v�>�0�c*p/ZT�ʠ�w���,!і	jx��k7/���O#���ep��lDI����4��{�)��x�V��cJ��8�Ջ�Q�Ì{�p!s������LT�?���u�u��(���/��E
�������&���#�n���E�'s�x��K')���"C6��G�|Za�YcSܙ�G|��e�o���^4鰼�Ӳ{:la��^���I�����U��T*&��_״nQ�i�+�t��5��[��,�"�ag�7���䥹�^�wj��,�SDy� �m��L;m�g�R���np���k�n�����e�Tw�9Å8�A�C�N�^�S"��PぃMt�ӿ�x� �[W<U_�!C�#D�\`/1�Y(�H-��v�j����ă"����s���>�Z��h�,_�th���Q'x/�d�_���s����a�8�H]..���XB괼Po�k�o6�Y�:}��fʻ���V�����܄W_��8�j�^�I�Ql~�1(�[9��{o�dy
�f'��O����ˬ�����K&N��LF<w�y(H�tī1�ީ�f����r��K��jT�������}�~�m��x�sԦ�I��z<W;�
���s�!-tqg���n�Ra�;β��XD�-3{���z}�*���G�X�qj�1lz�A�s]1	�hn�Y��cfm�La����%O��b��]|4���4t@�"�rK`@�|�R}��fn[��)�I'�/��(GO��7�̬`Q��k��|�nmҠ?�R;���k�����Ŗ��I��2S$������[:OlۆOc�V$�h���j�K,E�FC���6LI��v����[gw���x�Z�8����x������.��F�v��pm
zR%5*,©����'`Ѧ�}�WՓ�T;;��MБK�[�cOl�s���7���c��Կu
g&W��U #���ʀ�,��4|d�,`�e�K%�]�u�cG�Be!�(��7
��J���f���'�����Bd���[�Uq�R��j� ��>���_$������hW��ȍ�6��3k���Dr[/R��J���˔}Ϟ�K�LO
�<���w��-ԏ1>�=1j�.)��R��g���}�v`W���)�	�H��X������k��������(W7hJ���q>���� S���-�3j���	� :��/i���f;Ѓ�'Y�)��9�s�S��hт��k�@oJ��;����&�E:Uӎ %dL-��D�ǩ"�ܛ�]VY�Wcv�k�N#��}�+3;�V�,Y�a�9Ћ]������F�n��ϥ�Tf���z��0�|�$w|�
�3/Ap�?a\��H6�h������y�d�ӝy�������]<�2���k�J�^}�I������Trgӵ}���E���xU=,o<��_q�|_A�X�-�v6��Q���f�����n�(��ƌ]�\�L7�{E�����uqM�6oS��"�D�10
�Y;�ZxxY&	�,��؋�D��� �ۘq �����7|@EF�K��<�x@�	ka���ٽ��-jDb.�6G�jR}! �o�K��6~�2�S1U��Y��1��!��*qa~h��k%f��T4�I��� �=,?��5���72*WX�c��~~ �H{�Zs�i[� ŧ��(n�7��+p�R^�J��5��������nG�G�a^!���oJ�\!wx�����bn���J/��yw�i�O֡R�_��_��ɦ2�r�WyE)���!8���g{��� �����B�ZbE�6���P�n;��Y>9��#囸TSzx�}��)��J.=��� �Q<EG0�*l�p�a�J�1�ځ�Y��N�;Sr8�����
��6���2L']W�u�.��"�O���m^�)��`W4��Qɭ��Hx��=0�%�3\;�O���^{����s4��i�ҽ;�nK��-��|_�v��^��9�
cHt��؅��o�bbtBS�F��9��^�(�?�'	^`��$K�%�_�'��^B@r�U>4��a/�y�����;������pw�S�����jkkC���k��D��h��1��rE�Du�gM�=Ju�%������M�X��>LD\3�E�f��d�.
�$�ӅQr ��9�a@�,��ö���_�ƸZ({*��r	tW �M�M�*T��)(ρ��ûn|i2b$� ������Ī�Z)�?��}S���M��t{`
��4�%0#|�E"���/��Mr	���l�z�2�6?�*W���rG��O�J�`��A�g߈�H��jb�*��c�6V�߅�'��%���OD��x���'��6W���߻1u��0�&�z����	nL�V�uE@�}�Wp;}A
V̜�pkΰ��͓م�.�0tuqr(�|3P���Ԟu�x�N�Ո�MH��n���?]�f+�>C�a4.��n`�(��N;O��?f�,��"}�_F48���PB-��Yy�= ��v���k�`������A\_]����Kyo8����($��j瀑i@���պ%�F���{?V�^ϊ>Z�=�~�O�.�����3�?Ф�Qwh�􈐍�gd�`s�ю��5�����q����d���&����t�M��6��D�q�R��zҼ��uX��H�	y�p�����$�JI�]�櫔��d�$�^W�:���p)_ I�\�: {x�?+�\����I:�u:��cv眮�\-�E��O�SBq@
�õ#:�e?P�L�N�bd��S�>��o�-V�jߪxϣ���D��5�ܛ� ��:���0K�B��f?��s���<\�	秪Ly�� [#&з"�a@wJ	��;A+T��qm�&x�f1�Aʽ4�P�e�o�ӿ��؀�|��Y�1�T���t����X��Dt�7@�9x�r];��<�����,o��͍���P�3�����,K��ٗ�6]�Tv����v/AA��2�Y�N�1���Q^2hy����_:$p]xQ�L��~�-tl�UG�u�ݳ��R�dL��s�uCP5�R,EG�8G^M��V���_�CH��p�tŌ�>���ܼ-cs�c��|S��i��^�)��⻾��(#�9� �nYB��?)�O�Q	U@#E{��	5��y�	?�R��`I�
�@l1���7�4�0r�Z�i�. �l3�yW���_��E��]�c��$:���?�e�ˏ�B:}[J�a���c��K���Ҙ���� np���Ư�s(e�$r�4����h��Ix���-e5:O��ބܲ��qeb?ڵ�V�9w
q$��4����H�TU�MX ���<(���?��6�¥��9:�BX����Qx�?�"ؔ���}���Y1s�b!�m��"�p���Gt��l��a����Ūs���G}T���Ap�2a�+pno{��Y�Q'$�߲��$��V��o�}�Y�ga)y������AwTbIڑ ���P��ҡ��b�ɱ1|A�ģ�"�X�7矤�MI.�Z異������bv]��/�6�������F�g4��].�l�c{����gie^I�}��!]�-
d�j���64Ÿ��.��f�AtH����K��գ%s*Y;㤓�t'�0���Mt�ɒ����;u�_�}�,b	�AaWuZf&�2�>����9����ؗ�!ɢF�'uyB��v�&i��.�L���>'z���FOJ5N�E}i(���v�9�_yV��6����������ɗ�Kf�Υ6j%�s'�+F`wn��ݜS��!�W�\�����4/-*�r=�6%{��Z��J�Z ��B��E[�l�\7m�qߠ��u=�t|���h�{o�FZ�[�m��B#t]4>�zևd�ď��$��R��o��=.tkc�X{@�h��"<��+�W!�ǅP�O{$�Y�8<�^���L6:'�5��yi!1�t+:�K�sÌ��f��-���P�>��c�M�߃��$=O���ͥ���0�����qmآM�ͩ��
��e9�Q2�Tf�v�<@��HJ7�-�=8�Gr>����Rΰ�Lѷc�����R\n����`�U�_\�0}��|�h�Zv�C�����'+�.��)T�����hZ65��������|i(�|�g�yv8OS'=�e?*d�������h8�#�"���QF],I
��	����gK}4ý2;O�r��-�.h�e"����'C��r��=ϞhEy�;Q ��=`�q���c���[�r��2�f�bO����>��Nk�L� ;ӂU�n�n	z����h�~թ�ʧ�vF;?'0�[,���u=�x<�#̑ ��Hy;�����+���s�Z����E�%gȈ�o1U�����)����T
%�נ
iHlk�w�~&棝�o���V����Z��WeH(�'>I��d����]83o��n���\x�ms���l��4�P�L�~����=���`�c����������
U�����lB��#� �+>�PI,W���b몮9�f�L���J�Q�3���u>Y���8�x#${��=OL)Ϛ�O�Ӻ��XQH�9F�Nu(��~���e
�'v�~�����x2��H��t_��aaq��]b:�!h¤�1�-�T��:�0P^�A H(�3�<�N5�������k�V���GS%��k@�f'���E+�[�����@���t�H��EM�F�o����C��Irx�T��F�BIo��>�o��ݷA�@�&����n�u\?�G�M/Q�5]R�q�+:��➥
�*�f��젹m��,�Q�״ �:2�Sb��[��<�*B~Y\5�SWW)^_O�2�A4�xS�'�l��׶_
GgQ��c���R�\�a����;���x�������Oi��<���Dv��դɝ�j����>;�V�gg<�E�(��N����'������1<G�=���~�-� |,#���Zf�wS��戅�6�:֔S�Q�e`6��[��&Z*U�'u��J��eiY��wy �%Ԫo���`f�;�EXG�40-��nR$� Ě�cy��;��y)6Yk�m�(Ihm2`�"5�<��:���O�~�o������d�S�ضM�C�o_�ˉ��0��]3J�dN��liB�ï|�E�����{Ո�(s>fx\����t�=����?I��ņ)'�Df��mpn�8	�6���%#d}ux���M�/��m�⧶�ƢQ)�5���{R[͵�2�ZnR1	�zP�� 2u���;�3����v�D�W;��YmPǕ�$
�PS��T�}v�Q�N�h@#�Nvx�.#����d��<��x�̼̒G���.E!�x�p�1nRQF�Xc�!L��r}�ŧ�Z��=�&��FL�[n\��K�A_��Q��$���j�jEv�����Dd�����^�,&�L<��^]�H?��
(T�Rk]M���!�`%=�3zp��`�7�}�0�}�@sp��)b��k���]s��>��dn�N������� -r���k�}TX댬��rl���]=��S����ɗ�m�6P�%w��;p�x�U�{�yiл��5�S	�ǸLy���Im�w\B4�Az��VjsӞ�b�W�s����Jԅ<�!d1�n)��߸>���E���Ns�b����0_U��'�SyY�5�=��d��DG��1M����Dn�{P�T�*̄��B4-,?p������"\X����V������;��F��P�g�ws�>�fF�&:i> oM/����!i����.i
6�����@�FR�e|7nw��8�? T�o*�m2Q>(��mWj��R�>8�f�U(Ga}��rR��h��>Sħ�.O���������v�[�9'�9}0v3��_:�~UB���L�L�~7��6AA�u������U�a�F�#��kr3��],����e�>g��>i`�փ�篮��� �}\�c16�d9��t�3�笵���	���=ń�q�7��J��ג����I頠����_��'=(��z~��"bAm�Xx����r	��d�ڠ���8煂?�V�۫X�Gj%u�.LSBq-�����.wKN�8D�v� �Or�{���Y�����B2�Hj�����=�E���4��}�b��Z}>Z�r�$���JW,�U1�s�貗�.{����s���Xl$:|0���ً%�˭8c�9_#AϹ�{�F�e�^���.6��"��G�F�t�@;�k	��T&�#WG4:�����"ٖ��p�X�'j�]<���A�,�(����i���������[���%If�U��ͮ���f�ϻP<�52#���i�l �na��ף�IE�	�m��C_HY��J��1�*�Bo������j���R-0�Ds�c�G��־-�@V�|&C�UX����G�x�I�Ck�3ތQ��h��v#��;�'|`I��B���h��i Y���+�ٞ�Q\C����3q����u�?F�%�"����$]���=��V$f#\=)�`�X�V¨�ٻ��5�|�w956�Ȅ�`7_�Π�����I
G2O�!t��p��9�4�V�~��:��B�?c�S{��'�ֆd��Dl�ݽc�!x�1�#?�Ri���0��?��Ц�n�T?��5<���4Z89�=�I�>|��ҧL�;��W�#�LĒ�O�f7g٫lK�]����e�Σ��#��B�5��9��O֓���Ȋ���Mu�w�:_�O@c$x��H�+�Yx�BC���ћ�����]�cx�h�]I��۷������V�tl�\��ڈ7���^�MC����\d�I��'~� QM)4dI�c/��VwP��D��
���I��`.de���Se��6W[��¤� b����������x��e5�m(HO/�B�t�{,������睹�=�vh��)ʰ j��V�If|����A# ?s�myQ�
r��#5�縴�V%�۰�#��b�E��M7k�L,��C,�\�}���m���9��cG՘>�<�7EaĀ��=�#���td�܇vP��)���
��8]� $��4M�j)Қu�|{A�0�|����{q�xw$'A�I��V�Z���3ځ��ķ���5�\ ���#���	(L��u�zȓ���Gi/W�p��	�;%̷�r/Z�UXD�S~N`�D8s��=��֝+�iְ09�������7"�F]���[@spJ��ݵ�؛7�7Sx{s��/��V<=�߅hMv�����p/}����S��D�+�}�qo�j�{�K��(�OZ,��X��]a�F��
�xҋ�����U���ˉ���ݙ��P��o���s��.c������m�ז�OR���n�`Ǚ��ʒ�V'�O̊x��& %8�wT���[8��٧`�2��}���KO����W�xB��aM������mZ����b���n��ʏ'fx؞?���˩�فy��P̒�" ������V��K��g����49HkR�}��K�>��oeI^�ӟ��3��w��΅�QbM6�� �(8'~�
����?�p�8-ݵ|��I���W��\����Byq)��m��ZL�~��h�V!�u&��:?���S��U��mT��-�m�%�>2���q�{���ay{���(i���mU�?)<p�GJD�^���6B���Gq}��"���f{�%��Q����֔��ܣ��%Ɣ��d�o��_���U����2W84�t������&�� e������FrY��:�~����!�-?���ț�z��ހӯ C(�$t�H�}ͮ��D�c����)x�5[l�!� ��l�z� 1����i�p@�ݛrQ?J��v�z<P��ݵ̓N�� }m���{�nyR������8�S$?!]��*��s���B T�\�0�X�%o٦ �wH5cws���� �ۢ�d.xY��fSA��5`��)w�ˣ؜&Xk��u���@�d[�Z����Vo1lH�B��s��θ�\DH�K!�����s�C�?R$*b���s �
'��b���nj��tK|���x~N%MU��ѠwJ�GNH��Z�cb�,N"�]���V^zw��>��e���<��<�q��� f���Ĕ!� ���1�9�fm�\ҷ��
�H���h]K��=0h�2.��������U-,��m�·�0��_�×Y`���
N�JVU���&�p�o��a�r��e�%1����sϖ�KW��݊�
w?77!2��ZX����]�2��Pd.����\����\s����j�ۥe�� 5��%`MO��;��!�����h���T?{�)L��ع��! .i8����sي���{�/O�%S�N�i��}85�>����\�*�\%M,g�C�K�����j�ɫ�V����]?�(���ޥ0|W? �djfk��e�W���Ѝ�ڛ����ަ?�|:촆������?�1�t@�Mo�%����r��F��txd��L��-jࡅ�l�w�6#]��E
���M�)[&Q�Yi�Re��r����ʇ��g4�=��G�c�Ъ�:{�����y�m�+A&ny��k�V=C���^����o���D0���mv�2��5�6}�;ö�Ò�Ъ�����/�a�:�r0'|�F�B����'���<rR�8�(�(�"��JP�8��:�b=�	%,�[q���9\a��9_��csY���jqأ��H�>6P����P`D&q�bTP��'���`x�{�E����9^r����k=*ԓ��Mh'P]l1���?�F�V��W�����/s� D|�:~�5��#���dKo�p�$h*9�E��SJ �G<��֟��v�?.�1hZ��ק�Gh��>x������.������"�2n�ڭ�E��)���i\!"Ӽ����o�?D��nw�����Af3�|�c�u;y�e�����8�|��嬊���.�%��-&��_Fr���:2{�Y���^߈�[+�D==�:$�����E�Q�Q*׸O)�-��l�U��c�8�=Q����4��V����2��/]��\':��:���UBꔔ��:IT#����ۿ�v�B���5�ɺ�Kͷ��D
�I�U�z%i�`�Xb�3�����N��׆�pG�m�ECVs��'c�z��g�W� &�̆�>j�J�q>�Nt��l��+&�ak�s`K˺0��M����u���\�4z]]��i�,O��_;"{)�=l+��'n&���M�>�=�w�V#�G�^������Z���^��>��F��8b�t�΀���p�a�Ɖ1p�ɡ/�ItG������)���j�A/s@������BI͑:5>��
��/���jcĨ����UKd6>S֑򽴦:_"H�μ��r0p�2f��}��5�y����qL�g`¶9q�[qۦ�3=�yi:p�&m ��(�A7�PֵZ^'�#u,��*V�I��Nu&#)���q�@�\���.m ��dK��l��q�4�.����e�H�B���~������A�F�&h��B=�k�۩����J�>��KH���%��P�s\�z������5$
^SФ��+K� ��X/C~8D'��K		�d�˹DT��+A��{�a���~_��C���V��ǉ?���&��C���`��k�~^�6�ծ�:���6"��+'��.�œ�W�壄�����s�Z�W����s��bҹb����a�ɩ�)�	 ����oi���_E/�97�Y!T?�-��\�څ�\)2�Α7���v-P������.��6���-Yh�w3:�z�Y������J���u<�UM�6�1P�y2����	[=��²�Q��N_�k�n�@4�1�x�%'*l�'l�M����á�
�r��b� g����1��L��H�r��%��|ɨ���ϣ#�����z�:��?a�y�MT�f�4����_�[��Iذ�w����W���]���Jlo�1���Y�_^��Ul��Cͻ�103�ڴM�iO-:���9�_y�b8�m�\�~�
�s-41�Ȍ��|�z5� �cKGxJ4��S,��Ѿ^"��,�gXұ�K�r�4ť.����ڳ�ڧK�'I~�y����:8���P��.@u{����s0�ݮ�^�f�0]a+�������o��Qڙ����XIX���9�S���:��HH��r�n4�DQ�e\�9�+�zv��r�IN62]����`�0W�)��` i p�j���x��$h�يսB�F-2S��;,kC��ƶ�'�t��cA4)�nO;h�>!1A��k�EHBg���Є׊W�`�SF��Ͳ��'ispO��j�*�ت������8+���I&h�^�GY��9ox���L��и�~����'WH�vä?����8<� *�c�2�v"�Ư�`���&��O��S��C��6�N��s�n�'@PGz^ؿ��I|t�^pi�G*옰��i�V��<5B��?!e�Q+������Z��^0���<�c�IQ� �(�&�f�+�<b��	�Q��ɑq2�:�MN($����w���=P7�
���l�dPոv��X���v>t`����Wq�������0�xZB��mqm��Z�/\�N4�h�x�VJ��G�]R֗Hq��C���ɬ=:�)e������@�كu�1Y�$�����ݘ*X1���R�&��M�99�Nz*GW��<�*L��x(ڃ��ࠃ2�s�4=n��'�y�)�r�3'��5�#.[�)`*��QAZL�6GO��HEW���֓C��¢��Y0�6�/���C�h�-q�JW½��҈�]�rJ`g��wRp��v��2��>�-�s�q����M�����t}�v�!�ĻM�RDd8��PO̢��o��(�[��Gɚ���(�qj$w9�Q���-z�x��&���v�8���QǙ�<Z�?Fe=��8�	����_d{E\�t�=�B-阆f4�͹s�s���_s�����(�Oׂ�pQ�NN!W|*��t��*}��d�Ȟ��4ȱ�������MĀQ��^A\�0���.k?1I��+��̫�}��5o���[m�tEb�A00M�+A5�߃�{�{��P��9�hI��s�p��:=e8��N�Z�b�QB:W��w�y�g�:Y���ΓO�<���n_T3���f\�*x��B�N?��U��lKo�m��/��ۣ���n�/�Y3�5����O{QA3�ۥ=�!�Sx�����k�8��/V����dF�`�7sO$|��F2�Y�'9_�Dsgț*'+����'<�����+�]�*%�#N}&�2�h�&$��j.�6,b%��Ą��a6���������piw�߾�t5��՚/�s�� ����J
�|���;R�٦d�b�Ԯ�T�ڂ��(���|N�)5�=9uŰ)^�Jm�U�$���������2n�q�_r���(V�_�" [�H��8eG���\��š��S=l�7���� ���mV�*��jf�s��7p~[��r���a�Q��)����������~����3m�v�����\��xY(��+$�Տ��奩eo���W@P)�L����,`�5!�:�P����Q���L��}z�d��ܡ�N�*{"M���^���2��/�M� bˀQ(I�Ϗ$���!0&w�SU��R������3+���L����v�Q�|'�}�n�H�P��j]�?՘�V�Ŷ�&��dRĨ��o���;�~g�'�;,��`C�v#0h}|l�|�g��쇨����
P���:Y��VS,���.��Q/˾�(�K��J۔ʾ�θ�=�QMZ�k$���6�+�B��jB��.�L�9�7�ނ���8���8�d~�g�&�'�������  ĩ�ocW��aMtsq7qI���E7���'��[�-)�Q莘OHޟesЅD�(��W����1�@W�MqLPInE:��H�Z���Oa!��\���S���y�B�ॿv�P;Vܜ[�m�2r�[�/����F�'W��/n�5,�g������H?����Bx�Z�rL��[����h����g�ìA#M��9%nS ŉL�K2���lc|�"��v|�����Z;%��
��
 �o���B���f-��o�l�^�.]බ����ѽԕ���6�h�ڏD=HS� �z����ۅ,)�<#f�yo���Q���ζ��7�|cwQ���IGm!R]����Gr�.���a��Q�;�;I�Z�{N�E(�H4aV<�׍���WTS-q���Q?���7�ʓQB�F��4��/\Qu0����؋<�Ni�Z���BN�ܸi�2=Otl�-�c(Dʁ�m�c&��X$���_<X�t��Yo@�u�?��-�.��"�̳��R�K��V.D�_�4����� ��+��9a�1��ϣ�L��j����؅�1a�t+�����F,Մ�r�wO0�e�_n��qO]u>xޢzk^{���aA���a�M��Ҁ����w�IZ�� F��fC�N�{��w��c���c�OV9�4B���͡g�ؼ�������Ow��×��Ω_����B2M؆�3n��W#h��}�����l���uX��U=���8���,s٢P��%�G��9�� ��+u}�jSj1��qD�|��x0��.)��B��l�-�'F��|f�x�L�7o ���4h������ȉ����R� 	z�)��&c�k�\@�8HΨ|@#�e5�H����uы��R�erh� ��̃:���,�s��>B����-.Z͙��8P�Fh
J�]�
7�S �/���)�W��v�~�1�e �9A�[���6bSH�]45��qo,���wJ�P� ;{���`V�}r�W<��"���"��p%�]q0�&�X�����/+ �*����{@t?
�"ͳ��]Ќ�p:��1��呸pH R��n$�E���Q�����̉U�֯x�9[ſdD�0�r)�۳tʂ@�>H�.98�]�s��,.m)5����??[ȝ�b�w��,iI��l>L_���@R���#��V��%���('� �G��w�H����]�k�+�=�
?�nD�@0ǀ�����9�9<�2|���Yd�i+ Jϲt��5���I�laj��ʗ�e��p�����)��05 b��&Je ���g�?�r���ڀl�;�ُ���A��k��x�J���Y�^�9�Z�~^�4G����q�#����9JsN٩^`��k���c��Ɋ�H[d�4T���w�(��5�#���$y�8�e��6�P�"�p�����ٮgD.g�H������/�be]F��{�&&�Uk�H���*˔�H"�p���)�<2P1�����CB���|f��q�4���Xr3X��<զt�?XG&�\q����H�'V@Ց9x2<�HE�����o�q�*G�+�v��*���2-<���[5����^��+���W������X����Zg��������lB&:36�|@�)-��*
�P���B��k����!up\?FT�"�Q7δ��a!�j��дا��~P��(C�0ZM44� ���m���o��XHlC��;L��=xܲ������)#�l� ���:UFB<��$]4Y����m��a+,��z��JG�og���c����VZ�3]�[�� �DZp#�Wd�9+�bN!�;��Jx��Ed�yRt��lQ>��WY+V�h.N���J���`���<�2?����S��Ax�C����]R">{(�Ԝh���o��.�g�I�2;2?�wk�re��L�~�d��ƟH |����<�'�<�a)�o3�K#PAG�Л��r�X��i�*HtԈh�nh+Csa�N;k;[%&P�2Z��t�3��_�#���6f��#�y�2NkyPV��21�̀�V��Z�����Qq��Ʒ�q%��b٪(����	�o,�:a��IM�Ǡb+�:��GGba�C�ob��3|����X��a�2�tZq�9rGmW��(��C����r��[Ct����T)݂@{��z�MÈp��;�fb�Z����ƥ�Rr��~����ޚ@'�IX|�(e�,)���\�Y���}jDg�u6��Ҍh0���<��d�s���yÖ1��y��0 <���A�u`��	�GV�����47R>�c���#���ڤ?�[k��$�
��W�HJuT�=t���J�[]�5b��9[���CqB�G�ҳ�>/;6��O�w�%���`��ٽ��GC�Y����
O�`�`9��4��2�s\��JcC-u��dKS�c95"�|��pa�a�QQD>���6�W-�G�w�e��S p����:�f
��s��X�RD��l��sT4�55S>;f�X��}����� j�x�AG��?t�dEE�A���:	& 1A�x��h�h�����0��*h>�#�^,7����y�ꓬ=u�<�ֳ��B�����ѐG��Qp_"�Pb�
��\��$�;T�>��D���^0�|��y��G>�����	��ES	��b�55fߊ��lH�7���t���,�*���a�0� -�ޒ�̺+��/?KK]G7���d���fj�<CPH8Y��p�ͽ���_[�|���Y�0��
�4ι��
�fW_qm��YW+�[ ��k'�;��Y`�"��:�7o��T^
}�K'�w���;�Ga�vc@��t��b>��R��ד���b���u�a��j.����>��K�
�;Yy�B�I�U���/l����y(�����`�s@�
�ԕA����7|@7�kC�pn��dI
�07x��c�]�5�kĪ_y�_�-�^?��q %f^�6{�xƻt��(�ރ�:��qy1��\�����ɏ��0�EC�Nl�O�����������Hx瓶M��`��^�����]��4�s+�{��N�C��ǆ���0��h�J�'�&e#�`�K��g�#��ɫ$��L�/�y窑W^n��8Qx�+9UA��K��[ �SB��Գ׊��9K��2��� ���Z|,y:� ��k]�
:���ȣ��=�����j.۬ݎӴ��Rz<�p-"��q
~���B��U�ɲ�Nb�IN����*8�*6��9�T�_Q֎�
W��X��|^�wxm3q���<���WT7����;ɳB�����ǲϞb)x�clb�k�lve���2upsZ���	�o3L�� �e�}��8<�
4N*Mk�r��[��^��FB�	7 W� ���b�H�ށ���_���%n,�����mE:V��H[8��>w�û܃��ج�xؖ�6c�-s*Jo�_3��hr �����v|S���-�`F��y�x@�7��2����N\7��^�ݠJ��U3P.�~µ��X����A��4[�\��d-�M��L9���=����x{��!}l�����)a��g��^�	�}��f���яd�K���d�@�O�7Y�]����|�N�qD����Ȕ�Or���x���w朲�5���݅�\AT��N�T���[�'���2�E��:%ֺ=k�!7@T.��L��Vv����gݞ٥� �Np?O1�%c.�b���2Щ���DK�X�gt���֕�{ߝ�nL$@c�c/i�/��9�� +}
'�tM���d�p���$�C�c4�WL*(��dh��B�s Yp������eT���+�g˩�# ��w[����.	�^j�^��a��o�s�c?��f'�okeי@�ٖ�?�u��YD��k �R�p�`����F�M���j������d�Ѽ�@F]���5o@�bc��ۤn���;8���f(�h'�&��SGܼ*g�EI�T�ӓ\�p�����yI�p�\�R�?�
�('
M�����ŅCE�����ٟ�te��/��@��T��2�'퐤���&,�M��5-��K�w����R��D�y��TM�>0\���M?��!�/@��.���T���ą�
 +Rȿ	��=�Tܝi���1\9�yT����)e �&#�{�NZ��G���U��/��*~vLJ�/E~�MfX��4�+k�z=E+�R>�|�X�fwƧ�"��[�7�/R��|����!ڂ�(GG�C!'B��e[��on$�<e@��IRpD�W(ӅpjA0�$N��`W�ZB"*`Cs��:#��H��S������:ї`���_D�L\�D�j�M9����D@�$ǹq2BK�=vr�W>!ùgެ�+ŏ�qkz_��vq��y�s��5aR��E;�B�8\Z(6���.��s	���	G�N����˕�pϗ(1�u�?_���H'	Z1w�:�=����'e�´cH6?�W|�9�]T�)(/� ~I��F�+�X�����.|xY�/���a���s5��sxf�7�K1s&NX�J�\��)�;+7�I�a��5�=��?�|��׹;#q��~?�O�1�D
����`4���>h"�G򪞎���6dc硟�pw:s�V�������A=ʪ!�v�BL��~�N2Ua�B.N]��ǳ��8�u>� Hb�ﰳ:.��b��y<G�V`��z,�+��<�^}q`��څ���P�q餄+��(�W@	���[�f]Pnʦ\d�`�	�(�_����������1/nก���o�?>����pD�	:6��	��9��e����?3"(����!&�|p/^jc8���R���ø�k{̋�O�YU1�9Zp�I����/��,�����K~���m��S�N�c��9WUٶ�!���W�(&N\]'C{8�_�w2����n%/�6��Au+�*�n5PC�Պ�⟆ ��f��g�uP$l�ึ�W������*��*�3��k��ҕ�튄q�� �xO�9;�� z��:��
���!M\O����Cpq]4�!�N޴h�-b�h�P)Q���L;nA?>Ugb�Eשּ0���\V����j/W�N�u��D҈ �Я1(�_F^Ʊ�1��0d�N���ˆ眔h?C	���gk���ý�w�?Nh`�$.0��[EtW�7l�6����?�.V�&�J-��fI`BbT��U���Vu9"���)#Z+�|=���%i�r�
�:=F��|�h����H ��]q((���v�2PN�_��nI��,�W %K�hB<"��#�Pc�Ց�##�X��k >K�=�.����)�W�	����J�����;LG�y�0�U)xb���f}���0h�����
+���SA��M�R����3��
�WX�	
�<n�xZ#
��π�۫���y��|��5���G��n+�O]fNF�p��~��ء���T�^�Qv�a.�ת~H�8k�s�M��v��
Û��Ɓ4��u�#\T�������"�+3V)��O�m;r����c,"�@��d�9� �5Hnc��h&Ƀ�4��e��_�K��`z�!?8� ���%kx��������O+AG��m�m�q'��,ۙ!!�ˑ�\�H�m��R&p��p��� � �el4�X��A7�GȫT{M��`a6�#]fʢ��G����rO������=:��@���|��R��Tsugj���)4-��c&�'�������⇅)I�u�ЊYO�2y�7�<���.��>z�c�D��`�{�V%�]�Ü���_C�1��ՙAؒ�P��e�mǞ��+$C�췭E��=��/���Nr����)!,�'����p𢻠s#��sS��7��)f"��J-�>(���S/�u�e�p�IOC���R]ty���EQ6H[�o���ʽR��(�&ۢ�I���T'{0ɡ~��p�i������{'�cw�B�rW���-SI��>�c�5hU��_Q��b׳��̓�}�^Ġ>t���"x�����VP����*��r���21 ���r�
q�]�FZL��-��d���]zp�3O�!��;��K�6����%[ ݯ��)�#N� �*_"o�z_�p��y��H��nm�\�s��
�%?�q_�t��Ǌ��'cu[N�G�[����rH/|�D��d- oqŭ_6a0���5�?��1��%8a�j�ˣ���"��oe���bf��5r�׬���G�7v�(VH��	o48�i�*��c���G$����uY�a��j?(��ei}J�U��#�&*1��Gb�����m3K��ϋ1�"�~X�߬a�!��6�p�����8��3�ݮ�B�Ah�E��1�x)�9�q�v�lh�t���`f�8��0���O�;9;�$�g+O8��z�]'�� '�9�s|?����	�����p�^��3�8Uݫ��[w��:k8)
�`|��U�0z�H'�XR#y��"�ݚ� �ĥ�M9L�vr�J����~$��6���'�'n�5q](�A��XR����׫����-����u_5������ʋ��5��0^�\?�M�nxl�Yl=���椱��:��]��̎u��E���a�ЍXMY�С�;�����ڦ�r�pR���Y��� Z4��9��S�vW��Q��,��0���x�9ܨh

�#)��Z�u]���X`yCG�%u�8%����S�.o����4b�Qlϋ�k�'��T�JNM]d�
����%o�1ŭ������H\�6g�p5��䊮4�;Z�M|��;�. ^Ɂ�~�O�.�z���n`AR��4�@.-�~~�����kq�ft(:b0X��F^�����$7n+9D�ݻ#3F�>��Y"�r�?P��-�m��@]DBy�>�-�1�3uG<ۇ8���_����x���NA�����D�N���GC�!<.Q���Oڕ�R�{~v�]��,��J�Mj}�(:h�E;�ƀ�݂V��D���G8Em^�=��j���脔~�)�ZӃQ��(�z+."@�j��n_L|�/�sm����h
W�\s�;Y[�����;��jTqj�$I���9�y|5��Y��%�C�?u ������1���8A;��S��锈�L���('ˀ��� 1�.:��W�EuV��tTCV1<[�������k��c�ɋ�����|:m#.s�8�|�U��_l6\K.�N����|S1�MxT�2g�Z镵�-#3��e1���g��2��Ff�i���,���ͻ�2������#��a�ݤ�O�5�[��.�jY�{��M��lZǼ*O�h�?�>6I�).���]9������ys��p��
N	[�o�P��8�D��jUW����������G�K�=�}�ı~�鎅�tEieq� ����]�+Z�i����O���f �w��Y��5��zZE��}���Ɩ�.;��Ed�J��Q�d�a��,4ݏhD����@F? ��L�A�Un0ɭ�����O*`��>��]�G�oLσ�.=$2�;V�(3P�t�3N�7c
x;6��cm���-�d�
o�ǰi�o���%�^؃P@�͉�����!QR�v�x�^�����8�����אW���:��U������N�;���B#3%����ӕ���Z�,���2�%9܇��OS��d_;��kb�&�i�����D2*����s�ӏhw���-D����"��m���A*o
����r�����=M1����U����R�,�
�Ub���4���ȼ�c�c���+̴��1�����_�`����fбr����e�^gAb=zF3�"M�W��Ў��zA51�z��ܽr�&�!�)��Tg��	o�����%Mᚖ��{�S`��c��1���^md퀮��\=*)Ri#����~���焖�lb(_f�j7��"�g����&��%A0�>����F��l�R���УC�[�����;v��d��L��@�f���
�Rǉ����*>7q	.VEI�@�2���8�F�EuFG��Ћ�L���z4H?p䁸������)�i����X��ǽ�\'`W%�F�Y-|�������0�mbR���F!�`��T���x,m@ �_� �b���1$1����hz�+�TN*��է6���ik�z*�\d�j��rJbZ3�P<'^�!�LV��\9��Sy�	I�{~���z����|È%�WqhBiM��d�b�;Q����9�LƐ�͈�k�%�{��C�.f���}���n����5A�Xt�g�N��M���Xa�ӝ�W=h��������\�~�8���7��i1:�%X7!�#���=�5�.7�:��Z����AK"�FƯ[y醮�J��*~��}jD�Zh;�+�yP��ODZ8=B{���H㮞�Ҡ;��I�y���܉�尥����������1ˀ�tu�D���9&U��7�O�������}��#�`V���/�&�ɔH�a�
��Hس����CۀӛxЬ��3V�������@���YZ��C��Y�uV�5���'P����Н4e���mU	��H�r����-��d�-ŧ���B�:��[�u7Y�x����K� ,ɼb��#���g�(#�m�5]��w\���WK�����ZS	�"���<���UV^Z������	��r��~ѺEw�� �`�:� ��p/�(�7�D*H��W�⭝�|a�z"��7PO��z����i�A�3���<�[�EXX�d��6���奲����K�ȷ����)�W\mukٝoc$sw��08`��7��d`�PT��C�]r���e���6D-r��o�6u���Ւ&�@p�)Q�#<]�^.���Y����g]Zl���{���g�Gr�Y��<�T�)i�.���?=Kb���PF=�k<$����0q=�;���8��r�m`���̻'�,�@���0j<2��Bx��>J����Ig�ܭ������;C��ޤ�\�(���ōy��Ŋ��V-���'���L���.8�Z��q��(q87 ����I9�A]xj�)㥬��Y�x_��n[	Se����6rV�2s�\�?���� �z��UN�$_�83Q�E{y�qqW.�����&Aɢ��_P�"���v�����E �_X�j=;i}QXM|�Ճ���o?����.J�$"u�,�d��~S�ĝx�}�-��I��u)s����8�8������R�t+��V0H�-��ZN` �;��7ԉ��z��9�K�P�:���3��wU�"��rΫrLX�גy�8���\+R�u��A��.r���!��,sI9$D�1R���NH�B[%<q��&�����U��c�ƮL]rS2<��Qw�6fZ�D��ϧh���W���p0�����P����.܀	f���W4;��%q?�z�W�]�����ؒYTԒ�	b��E�x��ۖ���a�D��wB4��&7��@1LB���_x�^�҂��m��ia���M g�(^�f���7j�J�d��@�_�BE��H�*�ă�}U��e1��Fu:;q�lO�.����jN�e����ޏ�����:��Z�C�M�zXz@���[� -+��Y��I��+H��f��o�(���0�M#�>:���iw]u�<��}�r�i�w��CŲ	/cq�!0��>'��>���^�t�!�f�M_�
�~�HxƂ�k�H��zSB�ƫ�:xl/��)��3���%H��(��G�Q�]yAb�]�i���Z����O���]�w�{3�$?O@׽._S��{@���V}��㪣 hH#e��W��ӁZ"�D&0��5TU�tBVw�K�z6ز���Ƹ�ε�0G�?�s"'|�o%�ɐ��L֭�����E֣��Ui�;X����OᇁX^p�Ѓ���R[����0[	b�X��yxe�J�S����\�,����2�����1m�� h�߸����#�e�#���_F��(f0���TiR�!�F��c�L �o�KU��c@<Ms�K]��(G��@��$��sj)嚮��UKȌ���{�ӻ�!-IS��G�Q�I󂠽ʑ��e����T�(20�tI�T}L�d�9#�<��e���'�(dk�'��W�F髉nU(��=H]�;��r�$�2O$��HM��-`�����Y�<S��AR�*�|�I�"5�|/C9
�ȉ�.���D4�����\��5��e$^���
�r�8�4�/,	�<�4D���U�Q�K>R¯��Z�)K�%3�a\Q�y���٧b�Mήݑ�x������4�.�G۱)��'�P����l��^:�������?�˧+� �߼�;|8r�
[��\R�IN*ş�'���[^�F���˙���䣰ⳇa�X�����t�.k��9�� �Q��:�M��`C�c4�T&�>>$r������ߖ���i�+9������<IY�0e5c��L��',�@oj������[»~�ua�z���U�Z��Kܯ[���|�|����ё�ٚ�v����k��(�t���%/u�/�v=�.�ȬE���ĕ9�y�62���-3�����$\.D�E�m^����O��7PK� a'*���� �?��o:��h�EM�����RR��X	޾Ib�����6���P z��YW����k�vVBu6o+����}}�!D�x,���MO_�03$$���h�8��a'N�]�N��fł�Yg�����ޤ鱃�ԫ��J���$���ެ�$���T_ϴ����$r�v�CT]��[&�F�v���y�ue�u�Odбk�F<j��v�`�B{��E��Q������Ǘ_�}��NBW�?Ҩ� ���s�����dw�%�®�(�vS_������צ��/>t*s�#�u��y!����AZr�j���un)�g0�@ǖ%0�s�A4�������|�Y	�q��Y����@����tx�Xc���-ߪ�۩��Ϧ��P�E��q� �(-��&���׵E�cF�J擅������n�����A�N7>�Hg$`S\ۓ'M���h��oQ甹
x="�ѰJcZ�8����V�_��?�����tު�.�+8����n�e��4�Pv���ZjV����q�v�*=\MD�k������")��{k%?��4=#�ȼp�S���,H_�,%�m��<��j���͈�4iʳ��r/,kn1X\&S�pm��Q���:�������Y.WLY:n G���� $C��^ʹ�?�I܂t,�H�Z���uq�\���f��E)�9f�mf$K|7�Rw�������.V> �	�藿�z��/�^��euR���>��S�j�E�O'��Oxk�H�����v�Y�<�Ώ����o�Q��xʚ��T>_7�Jn�U9C���F��!��Z�:�g����L� ��-�t���zi�d� JRn�I=vn��?�q�����o�n���?w���Y�y�h8�?ZV�T��sru孡�Y�4���Al�`��}/�4u�Mt�E�qJ� ��v B�#��>w]#n$:�ȸ���hE
�@W#6a��r�QC����I/br/t�4L��믝��Rǹ���%����ar���Ȫ�%2����,~���C)Πlz(Y�]c������,���Zt������T�êx8R�]WSKvmW(�7ώH���ɢkyJݴ됹�~�@�Q(��`�Q��`wt�_�>��)�S<I���v���>!2���j{>+Y�o���� f��:w��A4��ml��k @s�~��/�)P��;?�	�F7�3)6jGlT���R�w�]E���XY��IIv�2���RT�>���O�NͲ�b�);��������q2/#��p�P�������J���bG�nz�ə$�Ä�����_s��F�7c���1�<�	�Lө�[Y>8
�.���oJ@��}]$��S_��S�'7���0?s��'�!�?�ӓ�El�^~	�V�DT(���Z� _���@��U�zn������Ĝ\SXz(��2gQ>�q��!�P>�ު�q�8�� 
9e!��k�}�^p�m�9�4V �'�U}��ʺ�۬k��,U�z�G��SX��P�V1�_�$���H`���M%�DEG��Z݃T������,������(���@$�Z�Ym��aJ?��3�����ϬD�'ߥ��@�[ǽ%D�o���&ȁນU���8����v���R>�0�T���K|���Wה ��DH��L!�	4����G�C7c�3C�f��^��iu��E�lu��7=CBI���9!�����V#�R��<TH°����ե���|E Q\?qbQ�^����s7,yl@�t�;T��|���Wp7,��<�'&9�[u�.:v�2�4�ը@{h�� �	7SO�b�I���W�&8 ~���uՀC����WN��7�`Ԧ�נf���.�_����"�ױ�`�ۺ�$��6��dŨ�̷�>b��8UYZ({F����u��hA��Y��<᧟96���G����$�m��~a���Q3 �>=�įP_CJ���h��n����jY>R���(e�	�1�F��,P;�Hrk����Ҥ�P٘����b���l{��ߡ�ơ��Fu���9k��N79�X��ѯ�!�yt��v��bI6��6��������J��˫�}Ҫ`��v��*�X�[�R=��ߝ8�I8�RE�6�d����c��_�)�V�f#"5	w�w"�2aS��n����Qz/AT/�D(e�"u=\7l���w WO�[p>�B�X�X���[�H�Sy9�%�{��%CHTto�Gu���0�yhW� �u������F����\�q�}����?	�]�r$�F�&K���p���	�:�$o{�d�+x�綆�1V� քf����w�;�� �1�V\bO4z�p�����[���nI�3�C�L34�n4��i*�@I
7Ax�� �
d���.o<ȏ��umvi����f����싄꼒l#���-���B���Y�b��VJh���3�_��d�_+��7�|�{�FԄ�U��̖�߹P(�p�H��6��i�Q>���w�= y�˷#��g8�����c�`�����д:0��"������B�n��+��e;��C}�a��v�ܺ�%�D�W�7����i#Õ�J�ˇ�Q�-�%E'2�F�)0*D����lq7�m<R��+����dF�OJ��j�{m�N����C;�o Icz�'8Y��g��7l\��H���?
~L1@(?�_J���I��_�Ub4�%1{V�Z�'I\񆁩l|#{�j�4�1ҸY:�xnǱv��>�j~Տ��VUi�nY�1�^�n\&��W����E�p`���L��Ak
m`�jI1�H�eɨ�=$D��,�������K��V���e�����S=���ާӺձn��R���D��e���v��@�+v�e��V �Tv5>N���l�ڤ��>	�x6'�U���q�#M���L�؃X��嫜N��]\&n���K-�/����[��l��lX�~fh����}�8�xR07|��]�Aq����9�O�2�!��==Q�N���O0��L7ƣB��^�5���1�-q���@���;>n�]���:�-o+��.72'.%��D@>�	 �`QQ����w����3N��%�-r�D�_!��(���'a�B�B���f������7%��z+R���K-�CHQ3��/*��ta�����-�l��J�H,�y��Q���dP":X1��������TR��E��X�B�,�u.P�Q��o"D+���L� �>�>QVq��ź�Yy����A4��=)�~b�H.ōߋ��j�of�#ᘚn��.��n��U?�!��S�@�̛�.�
����߀�}�hK��'���s����pjK�x����_	x��(�#{��=ʶ�{y� g~{���j5�î�G�bI����8�{z`���E9�'�Lɗ�bR�3c�S�6�U5FӅ���b��$k��[�֢�#]�??�3�}�XQRF�u�MG��G��"��;>����Ҙ��(FbI�,��s<�~�ӈ��Ʈ�M�����W!q�1�ڼ�E��z�Bt���a����7g�p��&.���5"E�M�픳Bw�m�_���/i��2��n�[壊����AI�F	����
��h�0�jΞ���Uhb�֕�WC������e��A�|4�z1]�,������I�5�r4C��u͇ N��^�".rb�q���C��ގ������;��ϊ�m{��KK�
�#t\r�e gI��W��N6��ca�i"I�{��Tr�zޔB"�~)�@P�l���s�\�F������ٔ�F4�W��]%��M�o��(7�K��u*݈�Y���]\,8ɚ��쪻��&b �a����j��^���ĸ��=�<(շ2���j�Z6�M2Z
�
vSm0��C�d(��W�?����3��_��BQOR�W�����I��d��ai{YMD�_�J��I!r�2ZKj���o�sƁS���x�2��2 �Ԃ�,��]�z`	����
�-�1�Һ��1������Ҁӏ\�ഹq"!�O%�`�u�F��F�}Ͽ�P�s
�G��=�=r-or@�{�����@�^V�W�غG��B��ҵ���&��s'	v'�2�5�<�&�l�a
uR��	��	K���@�J���8�3��q��:\��݅���Qc���@��"u�n[��W�Yn !��a&�Ӗ~2d\;��(�S3YO�I�{gy
�J	�!�}�[�B��ѧϠ2�U���q
"�'�=�p&�R�\wX��?�۞�4a�*�?h�X�;��ٰqu�6�H"�M���$>H�,����lX�YȪޟԔ���[��-���s��v�sie p\4^��D���5&��4D��mn�k>��ZqQ>w���髟�]V�c1_���30֧&�)娲
ϴ�P����BJJ:�l�%��s1�Iu�d_3�����8��_A���S���_ |�P��r6�Y�]�`c+��9�C4�<��g�w	u=@g�M��(���`&�8��`wy,3�=!�ɔ�l\�"ȍ��p��Czd�a8�ې��!7�Z�d�*^��f̯���+�xM��>?�ʣs(��B����2�P)�<t�������6��|��ZBJ+�V�S���(>�M\{� =%�2]8J�ȼ�ND��D@������d	_����]W����wk�I�[�D���4*��9��e P�;&N��y�����4H���-_��+�W_�o����A�Z&��ah�-j���
������6��.�.%E�2�Rk�Q�Լ��{�"�N�O�H��-�(4E����ӕW�P�LE�e|i$N8r�c�S��-f��):�3�H����e�<`���?$�����Y�Cp�u��SG?���~��mkoR�9U0����%�1��3�޲�
��ׁ]*yWXr�3����R�&�0Pw���]=KRP��>(q���ʋ�e��硎�篽!6�!�A۲�v���&N����@�[g���sWe��U@�ȸ4�R^
��kW�-"�I,�%��_+^�[u��<�Gx�D�� ���d���6�B�e �Q$c�C�`k	��@'���/c^�k*ˠ4��(O������ϐ�	?Ȗ0�Ng ٬)	q�Uw�M-�N�o�3|��%m!��\z�Y����>ȺđA� 3IY�&R�!&�!�n���PqUjT+{E�����ӽ0�i� A"��zl�^�k�tN� ����GrwX�4���L�����S������Uٳ�@OmP���a�M�鱺��D�>���`�ٚ���L�Aoϯ���P�ϠLNk;2��z2��Z�6�>n�p���^�^Y�(�L��[֨㳧%.���Z���Y���%@w�j��<E��M}�|ϱ�x���?ş�vܣ۴�t2O_�wV��i/�����f-�L19�FJ@���x�nρcR~�g ��)HT�7�AQԣA5��W1X3bĪ������arM y�bX���p*~���PM�'�
K3�̷��Z3L����4u��1�q4���?�X�Z�p|K�EMf�p%uAs.��{�r�?��YEY��>�F`Em�� ��\���Goۈ.�F�2�py<�r�Q9�+;��D�r3��Ќ�t򩎻��kE`��x��m�Ԉϒc�e�jV	C!xCX�xM�}��?�.���v����C��8�� 'z;����w�Nv�GЕ�N˺����:���m��ɵ�W`kI�7#T��7����X�U]�h�E����A��LxL,0�~���Sx��G)���IP����������.���~�+���`�*��f4�G�
�-�'������� 	۬ȅ��ȝ�Q<�BlT�ǴS8,�Im�g��!~��!7[Tx�>y7߅u�XL�;�;-��(|��v��eℤي��������0��o�2��j�VϺEЪ;1ٽ��@p˗?��XX�@T+C�o��J���� H[��l�M	����wKW �y#�*�Jt�T�K|�U+?A;=B�!�D��z�9�}Z�=�X��\7��Jx�g0���U�ڍ����j��n�kp-�f�7�]#�yYU�*�/7�[-�
y���Y�)�wi�.�_7�ʉ���ma+:�
�*��?)\��P�$3"Se��;��C���I����y��r���k�";�y$����B_���=dPQ>�൧�/#+ߔ��\4Bq�ęq�I�f�z����W���'5��v0�h��!P�X`|��?�,���%�,������wt��h����D���wꡈX���D0`̯�Y".�oY;=��}T=��)�ֲF����Q�:��
;0�%r�����[sj��詧]���a�Vߧ���_�]yM%�#�j�9��]0��k��Q�H�6n��~��wE5��XwRJ�$�k����fO���|�KĘ����F���Ej#�0���͐݃|�;ڤd��e~'�dXve*W�b�ʈ
#�)���K�R��~���w#�uV�	�>�ٹ�h�����j�Ył�<c
}�t	��/��k���Ei�p{>ԃ���W�T���A R��[��;@d��ll`x<���y7�� 7:YHiIY��h����(o��"�HV�+�� _�]�#3�������-��}"�*l�2�>L��� ��R�����Ʀ[]��M�BaZ`��BL�@�Օ�a||�c�Ќ���=|N�P�m��	�m7M�����8B��gڄIYÏ�k�sB?� zt%>��:B��u�TK/Npk��̸�J�+~�8��ڢă�]3Qj��%��� e���r��k��Y�=!4W�w�����~1���m껾�cy��UD���F��{8�q��_�9�� �X��9+���կ�����ܺ�2%�ǰ ��,���@��|�P2`Y�f����P��ʳ�9|B��{;9�/[�(����k�4�ɛ�P�ߺP��1k�a�?ߥy�{�sq�wی�ew�zeҀ��r�r0c�@Q�	�׉5O��4y��QB����I��fH6����,n4:�yz�	�z��!b�Ν�1]��e��8}���L�M~���=0��E�5��yڠeڧ[T�4y[)"Ĳg֚��ّDB���jk(�P�r�㮝�&��Wo ,���ч4��g���:�E��뎦�Q���M޺��<Dk�����nuU�7"���0�o����>1vz�����pYt�x��4-�s��R6�y��ᰔ}Oq���]-�Y�[�}�ҩ_l:�-��ORf'�Ee�����d�B�O�s(\|�2Bi��,!�Y� �|p i��(���P�@���IΏeĶ��(�� �Ͱ�c1��l�]Pڽդ]�
�q�^�6?����;����Wo�		�.��WZր��q|�ZY��N����	��\���6&���B��]>��arh�a�p��F�w�b Ʒ@:5��o�F!{��e�a��gV���޾�ģ��n���~O}񜃽�#��	�\.�d;˛�C�go���ӝ��z�Rש)�����C4C?�<��Q���*)D�N/�J��:rª���%.�>�aq"�rg����نGXC�
��7�wǦ�]�N��$|� �Y;�o��U,���
�5��"�K%�1�s�Wx��O{S-�nʊ�uut�e�����G.��|Tl6=l�߿����<K���@�5��������L��B;f�6���	1Ni8�D)*����⿊��,If�D}�e���oS�qr%�i�z��hO�a�fI��0�*��G�*�5C��0�5���n�־��t�C*<xs觉y� ���H�~��g� ж�[}�W<9�v���5C=�K���ա�d�3��ʟ��f�e����/My�p[��[lY2q@cW��&|z����7�*�ו���9�"��&�P�4��u�k�'�.��>��\P5a�����1� ���d�۠��t��vB(O;A�"'�[�<R'{YS��N��� 8�|��*��T�%�*�7�髍�`�ChNx�kM����|�?���6CFl5Q����k<�I��I�-�	����+����2�g�2�xJ��]��AT�$�w�T���rI�����������d�Gǖأ��R*�У��p���S�@7[y�|���LI/������TxSֺ����1;'��Q�-:�l�]A�v~����;�����q��P|�� )|aoE0�&�p�]!�waDWO%�+�@�*|���8��i�0ii1�l�*�R�q��G��u\�0���A۲Y���+�����{@���D�,]�� �#��?���N}3���źC���b�9���W���ه73��
_-;ꙮ�/��D�3#�+E=D�IBZv������,�Ƹ<o��2�����-����l Xm6 ��ة���A.���p)���g�(�hS��4.R<G���=E�#Y��Q
Aհb?�i��Zy�y�Z)FF�R.i�{7�yp���b(�#��,�7m
?q%$#�-����Fy��0B>�p.�a���9Zȫ�٧��m_ậȷ%�j���kۤ�=�URdD;���qH�)d��VD٘4G7��HޥQ�ݓ �����m���n��u��Ǜ�؟b_9:����dڼ� ܽ���s~�q6���)�u�ڀ���� �y�.�y�i��t��}�a�y(&2�;��7�����zYc��h��'�����:�|#��E!q�E䣢⛤ϵ��|��&f�\"�Qꜣ[iV�`���p���߆<L�Ň�5d��B���'9	�6�ױ+�wox�b��]	��J���{���m����l�kX��̈d5I����3.{�K�n�f��h�z޻���i���2
�e����y E":����ʎ���o�ʹ�dt�{W�;A�J��T�����	J�7x+M%������!�Hr,�Q�g��g��,Ա�=�gB���n�vI���+�=�<�
�6��O�d�M�!e"��%7��y����(C����ց7s�R?�r���#���ֹ�z&S��������"��L5�$@�3Y����wH.�j���,�3���JW�ZkӫX��_	�&[�k��k���ݰ7�v���W�����}�&�i�[��f"�|j)J�G]j��{��r�۞<M�����x�Ƽ��*w&�/	����޻z^8���
������x��*��e`�f���#"=���z�������WHv��a�D��#����ӳ� -l�w�g~�{��m'�c�|��J��ɯ�!�"_,h��[�|"$M� ��i+��A���b��:{yM�&8 2��1�Lj�<,���:{��V����Se����\1$��@:M�Q�~�o٩'��	ϖe,g8��ʉ�,��<�U�ɕ�kgu��XM/�Ⱥ�0�@Jwx��A[9�� Qv��ZӈD;���7.�F�iR�}��.+��E�4b�7���V����=%H$Ȯ��W�!��k*����n8�Q	�9��{������c:�K���G!iI+��x{M�� Eh��T$O+h8�@O�0mӝ�m����-����X�y[Z�JD������h,x@n x�"Ҝ��Zgo�����ѝ"���q��	^��-�{h�<��;��#r�����h����O�=g�}�_>#��N�~��t��j
3 �����Or���yP�ek�������^�ߊjb��OY��Jzz�/����&rL��YH���9�׸���޼/vS��٩H�M�{��b���ѡ-~���	�	O���8���=���]c�,!��#�m_+�k:As��M����A���'X���%tS��6� 39誒�lu��a}����n�8�X�J���!Ι�t�K�&�]��&?��-r�P���S8�9�ݸ�rqj|����ސ��n�D�t����З(������0ʍ*�Rr�M�7��㛚�C�74@0J=)Ŝa��<-��D����x$�����O;���[��G�`�To�_W�m	����g˸��%1�(��j�#B�h��k�3�:X��|��!E4g_Y�D���W�ʄ��(������Je[���e�|%�����6�A-	��}�Hl�΢=o��?��IG$4�L������7(ۥe�{;x��9�#[�}�/*��v�А�ʙ�K���c=���ˤ�v�����'���|���۪����?�=R����ڗ�0n/&k���@Kp]h��u��2ԦڈI	���D���.<��3��l��ޝ&�v:a�u�MO@�X2Å5le�~l�6��M��<�'�o� �:$��I�}�x�n���RC�G��h	q�"���Dl�\��d�Җً�Re}��$�<H���|[��F�@�b:��kE�]1.�����?XUȻc��3_/Z�ǞhW��8�� �qN"Y��������~�o�����+g쬱L3�Nh��Ì�?)M���[�����Qi	{'�����dk�z��s����Oi���~Q��ȼ�J�^iq��v��=�k�����k���E� ��\_U
_�L�V=Mgb�1-!������<��ɏa�y��Z!�Vo��^�.�K���6P��Q�����`Z~ggu��m�X�iD8��SG�YЊu�N��(?ޤ+�z��N>�Õ����m�n7py���<�'�!�H(�O����8`u��$͞����޽x� �,�Mx��aT���m�ό'N�:�پf�����l.����ر����1�v�L�뫛���x*T>[�B(��nw5/7JKAHR*�z��*�&��GN/���*�x�����8t��Lp�X{��2Eѻn���J� �j���0Ġ�5\1a�G� ��9�;[Q#�����Z����U�Y����}"�g�sg�Ad���?`�"F�Ε��񩎶���m��{ze��
u�;��3�����d9V�~����K^�Edr�Ӣ�X�I�Q�b�#-��[���q�81�ކ�#���Ԯ��L��.A�*$t}�23�@�$�7Hg�UJpZ�%ǝ�}� Gw��g�V���B��pL��x4�p��N�~^�������rm&��q�ܙ�[9pM�â�����^��8J�<u~���?t�ͽ]w�%�7�3 ?;�½z��E}��C�Q���/�m�e*��wr�G��C�����ݜ;��[lAe��N/��9���Im����X+��F�
�*ah������C"�9�*8΅�K�u-8�����k��@)�������q��-��ԓ;�"�&���f���p ]�ȓ���ĩ�t��o�s�aO��	���;� <��ٿ�\�S!5[7����ݢ�ԃ�>��E��\˪�����S��e垜E��Ϻo�$`A�]�c@�ڇ�@�hQ�/_TN�m:l.6�;���M)�����J�!� ��j�Pn[���?G���k��QX-��?��ݪ
$|��(+��v�K�ՒS:�~jm6�.5q��N�y��S�������Q�Z�[�E��d�Uȏ��f�����m�#�xV� ֳwg��Yb����޽0���7u�uÆ�̮*��:������e��D���Ǭ.؆V":��7q~@��w}z�;�?D;�ȩpB�q�i�Xݼ��fJ�b�A��|�����G�m}����D{�Wb���ɷ�[|+�xX�@[ 
��*��[t~Y�;9�D#�9��ʑLh�T*r��aI����}�je)q1�?���W.*�-A��I�~#������;	���T���ɤ-õ�e��ꪄ��JwĮ�W�,V�6aFzÀ�vdǾ�AW��e��+�ɂ,Q���]V�X���,��$�f�΃U@�~w���kψ@�O����H�zi�wK� �Dd1/����,1^�g$)v�u�{���A"JN��d=�j�`m�P�A��d�i��"���,?Z��-�l?�(�Q�Fij�?B2����(�hS�I�dl����T�wUDhM�co��/V6���Y�،-|%�$*8�g|4�@^8��;l�\���G��ٛ�]K1Q�����a`�p�Q��]{�žu�$���-yB2!Nj��d�
��.��.�$])�P<��F�e�0/�"�R�ݔؿ ���Y�_k��&��=eM���Ră��#��� k�����^� Q�8�9�P���'�����P���8L�ű���d�Vb�烙���4�(­�y[�5��83��o�!�]!}\�7��A�:"�g����$� ���^���8C{�p��:���N�!�N�3}́����C%f宔�P6�˻*~R�X:g��3]:��|����£v5ib/�+L�l=ͪL2r�,��!_Hw��X��޳d�B��O̻�l���[�s�)���⠍�#��
9F�o�<?2,��g�>���`�XE�=|HU펖��(�V�[G^>A���+��~�̰3���k�҉�fNVas���a��J˧"mW�^'���x���vXzչ���[� ��9-�����6`�ay,I�F9�sB��� ϐ	7%��Gb%�OZ%~r�tG��s���ir�]^�~.��&�r���Bz�H��E�vLj�C�ۛ�WEȱd��*fI>���O���|�[J�<(~��}�"��T�e�ފ�*٬i��SX5؁3�߸z~�r�V��/��ҝ;��
�h�(�~�JX&�E�Y��I
�)*u\=�A��aF8ͤ���5$���^kCȉ�G*�(�{>9#[L�e�-Z�l�(6c'auY,*Ѝ��-�_I�/�� H*D�r�:�#��s�F�K.Vd�E>ڑ��f�˜��@������ὦ:%bhJ���CJ��x�,d�򉲾]�P�qEJ�D����y]��Fb�� �I��D�Na�ۂP�Un���F6OEXʾ��o�x�����B4�7_"�e����E,��(44��8�PO��o~�fcnt����rfVI�2w�pCL�Hњ��hC�6��.��IRx
�sF8�6	����A�{p�%�w��<�g @�W����F�'�8ßɊ�V]�C����yK�GdV`�0N|R�f���;����$ë�I[�QP�;�&�fn��y�ㆍ��ϗ>�}��-���O}�d�k4r�G]?�ʜz��x�y��'P�\��Pe$�_c~}�R4>��g�I��->�D���l(, ՟	��E����͚N� '`\�	�[�>�tKy�V2��>��ۦ��%�
���;1kI�J~I�Q
�:�-��᠗�Q���dM=qb1ٞ�N���;{���Ë� �O���(?aUt��g�����h	ln�L�����%m��La%{<�Jr����H��g��*�%D$Va��\����]Wy���3|sD��C�";hOj�=g�>���V$�UFg{��#R��}c����o-��']��?�W�}I��i��:��E@���o5���бI�]�&�#t� �XY���Q�ne��^��O��C&�$	��e����O�p��<�|�l8m�6�V�?�4Uڵ�^��0I��WP�v�X�V���`屐h��d�x�m�����w������2�/b9,�4'���X�3�E�l9���# �������Bp>�p�=�Q�슣q��NX�ןY���To�U|?4E����v�8�z�`�Y�U]r5���:ҵ��WJQ��ɒ�7���3 ���P[�K�Wli.T�bJ���L�)|����ѵ|��9�Hbv��؞�-3��L%L�1&���R��hm%�<
ZwG����q�ew�ͺ�x�N�C'���(<Qf^D
M�J4�n� �Z>���ӇV�.s���VĒ|��-��W;E��;�8���ͺהc4���Py�����[������z��B׌j�";qk����
��j���c�\�2�}Y|m,!
�f��!�p��Ԫ;u�u�^v.mő�%�u����m��F��Z�.�v�J��9=�i�ۋ�5�BZ�>�)z9(C�-4(2yy�+�zG��]s#�<��_���w�[�R�X��^nY9�P����n�( v��H:�f��=�����Y8��	Z�G��4�:���=�+w�o��s�y��l����Ċ
��%�?���6~s�U+z�F������1YFY��,��o �A�e IT�7tw�A<9�;��'�K(�p��.�'�:1���ki_�[��DinT�'w��MJ�h��M�SA[�g����7~bhD6o�ooT\�<�`�����X�|�������0�����]䘉�ˏC�M���$�����}�@Ի2i�/�1�,n
ps��\��-�PE r��x�A���%�	!7_ ���� ڃ,[ȣ�_����C�s0��]l`v�G�x���#���,�g��g?,d���B��D���Z�O ��NeY"�ő�k��t�^�����l�,:�E�T������Ų�����p�JV���]Y�p7@�]�#P	��)+G9v������c#����V/i����s�΢�-{D^�I�`.��)3/DN�]�	6
���o�����($pu�p������(�'��Yj.[g���gR@������t� �m��}�vT�ʾ�k��2����3�ff(�%��D��z�ضu~�[�W�6���sq&^��H_��ﲚ�3"�LA/��m<��D~�(2��0`PJ��p�aIH�M��R�
Ӑ����Y���E�����- g�`�v?U��΅�fB�ǵb����n��(�qS;Т��I�|:ӍZ� �<�4�c��hc`�q�_<�p���β_M��]��\�۵��D�A�(E���e��jj�fTq`D��B�3��i�|�u�LrJ�(0��Wz#`5t�:�ٹg�������h���
��O�e�J7���u��j�%��	=@��&'��=��!���D4�;j�T���]�В��\?�V�B�Q�uΟh$�lG���}$z=�� �:�▸��M�mD�ͧ�'$*��Q\ )��z���Mjj(����������T��k��G�pH?�	l��n7�ȟb@��{?�Ќ@���nN�S��K�?�S�,���������Q�~�x��-鞾=2H��� x�hd8R��t;r�xQ{�O��=�7��T=/Bw{��J�&��0�K���E�'��@L�R'�������J�Yb��f*�����`Ʉ�E��oO����h�Fwuc��U�2<�ץ�8�f�My9\�v��xC�d�3(��8�`h�������놿Hv�?�2�=Pqh4׊�硧� �e|������
av��8�ކ<*^5���gpH���x����i��P�r�a�L�3=����6�_YM���r��[��K\Tg�������.�z7�S��g��Lr�8er�K����7�u� l��w�F(A�8n����0�p�)b.H^d�\�5hA�[�(����So�jSj�M�����c^�9l���A��
k��ƻՒH �Gm�d~Q��
N��4���+�|�r11�i�I��tTN	�F+SB������mΪ�����0��y{>x���=�N6�z�"~���t��rV'(7�7*�w���F��ue��� l��v_� ��$����WӖ���SM`�.~��U~/�$��y�&��O��f;>Ũ���3][@������KNt�d6 D�]�̎�q��A�[�������١��Kc"k<��a-d�%��O*��[�QU��E<32��0~�>fM\��~����[��0��)FwG����DA{�A/`I�B��Րiu�dJ%�#{&���_--��F�*���>��Zy?آD�X��5_\f�	�S]ոCW�LL�V��O,�oI> m7��WGM��^J��,AU�<;����h�k�PQ{t?U�h���#��9!27�_6�<�xD���\l�y���A3r��D���G��N��k���lv7�T��K%_�Ryg'V��h����ޤs4����]JƯ{@k��BB���*��ğ&=��,��Ou�0�	�� ���#������[v(GG@U����$ӆ*���&@.�>ÿ�`w'�772i�����k�ufye��ԯ�/� �c��]�e��|�ߥ8���EX���[g@6��V�Pp ߹x�N<����`��y���p�r�GjVNUͶ{4Ė��H%A�_Qe�!����UQ\ޮ�H��Ͳ���0ȫ�+]��b!�E��>b���C׌�v���p_x��^�[!�>W�1��ށ��ؕu����~oC|^N6ߖ	19�Y[${b	RW�12�J
R̇��}E�-�U�)��������A�����E��S�̮7?̸�,����P7����`l]�4�T���ƥ�15���'9��l�O�	%uD��a}E�>W�0^R�9*�6�4H�+��"bg(�|gʏ�O�oO
Ô%�ga�o���8A�B�Y���6��ϡUσ�su+9t��E�e���"��7PF⥴�{,S0լN����щr1j��K+���4�tܾv�&9�eA�dN7�S�Z�&	n��Y=Ո����Ĭ�8_��Op�U��ȕ0F{#bE6To��^��Z<��8�*�@a;L��BH�W�3^��Z!�㧙����6��bVV��<�A���N����ɝ���w
X�L���3Εv��?]f�yId���E�V�k�I#u��qU#�Q��	��0�v�F�ܳvx�Λ�`K����8�|�\qC�K�Bpq_Kh���edjz j���MV��ǻJ=YZ�S[��(�Kaٞ.�}���2�W׳���@�R��$�P?1��F���&���p}��4���MB4`W�<��ƾu.����h�����e��d�圔~,б��6E �r���P�x��=�4n���fC��o�+-�LZ�đ�đ��o���ϱY���'��e_��.ö���YK3R����0���,Bve�[R�p��tJ�����u��|����qL����!�!-{�S�K�@0�띚1�ߘ�ϡ;/% L^�"8:9ω��&���hA��S@4���B��@�2��;��B����{��[��x#�'�r-��Z>TŊp�Y�w[p)�L6(���iY��T?F2����V!ã�S�;c"��hy���E��e�lt�C�ՠl�fn� �/W�-�������"4�4v埂���zK��SO5��:d��oDQ����Y5��O��ӦIZ�prs!�;���L�|�|��P���=ʸ�(��CITy�4�\�"�ro*Q���� �8�Qa>t|���9�"<��7R��� #f��&�F����W��呏�U��m�M$�̢���٬	�A���L,'�SY~!�87�ʞm �6���e����e��2�����	9_�2/�:��J=��/�v)�Ԕ���� ��q..�lb��묓����5�ݝ��Sz�@�U1���2p7t�E�eс{�L���5��"�y��4tM��QV=���U��硑���3�9t��ʹ���ׄ��v�t�zX�q�Dр�9��r`��_*�f�<�j��C��Ѻ�kQ�+:�K'�m걒�Fc��~�HK��8��T4��Z�Å�G��m���$�~&���d�t��˶-:�M��⍞U'}̀f���ۇp3<��� �m����?�h:������z�7�\zѾ�bZf����e۹Lʱ-B��$R&AC��Z�w�M�b�E���]�/j������FS�,���[�-Հb�� r�d'��m��ʹ�����6�X���Մ�@K��t�����?�u�m�(�ʒ�ҹp_f�RQ�M���'�,���Ȑ�c����濤�Vrn�����:���M��a�]+%˭̩�q���2�μɐsxX���h�3Pam>C��}J�g3�j��ǰ��yМ7tV�pn��s�¾�E;%�
�+=�+S�Z�1����rʴ(Y���8( ������?�y&���ʝm��P/($�0d���UF��]K�9���Ȃ������&h��&_��:�N]����u� �����nPߑ�` ���N�?�q��Y����YInA��7���֞�V{�ԏ���NѬqw:<�~�s_���Y.�'HɾA�}ݳ򢃠ߨzo_A�%��kp���a�B�jбoT\M>�|���?x��b�HH��g�L�4��9�Rc��S�S��ӄ�L&���|_�(B���(�~pl������uJ�s�-�Psӻ����)0�STU�������4�ǒ�C��7:)-Jb\�8$�/�&� ��:��>�̐Q#)�	���3	v����~X�[m}�}��%�TP�7鹴a/u�hs����=��e��b)#�DQ��$
2�x!K*�����7?pԕ���X�GF��I��W~q:K*$�	��z~�'�	+N��-�oM�U/G�{O�I�4��Kլ]�Lj��  �х�J���OE��@�'+�{{�'o�ax_u���F;G���SY��G�����|�k
{��{_�K.��q�E0��{�u�G��&A��v�nʺ��0�`C}��t9��9XP��v��E��a�7:` ;��C�B�������D�&�9]\t�W���S�1l�������)���j�.���p��t|�em1�qc�}����Γ'
2���Y��)*ku4����궮~K����B���Hխ�h�QPj��,�܀jH빺��|�;Ad˾B���hV���q���=x��j�]��r<�Qc���Xe�s�G�ɮ,��ù&%��8f�|�DI7���P��ChیѢ�Ǯ4�x�]��`m�x�������lB{��Pj	�0��x�y.�+!Ѣ�1�����'K)� �hC 1�d߰��"�=��Oaw�g�D�1���?҈̅.R.Te-̍�5y8��P�F���Tɸ�V�Þ�4g��i&��C��iJ�9<��6��ߠ>��)�i��K=X_�/�0 �{���P�ή���XYA�[����#�Q�ؑbEt����É�탢���̈́�cڞ�B��8uɗ"C�x��Ϣ�7��
)�BM�#+����H�$vL ���uD�|�}�ᴫ3�Ԝ\�����j��D��\��&>CF���X�p�H�����?�z�U�(nlԆ���(��� s��i��/�7�S8��׹��_ϕu�2�,9>���w*r���>���:�Rj��r/H[:�� W�~��~Gq�b���M��!���u_�G�uŁ>>!�A�$�(�
���$0C@���?����M�˯o3�X��{`�O �w@�Ȇ��&(i�fL�5+�.pP��h�R{5NF>�}��P a��_ L� ]�����q�������XS(�N�W�{��هy�|�����4����G�Z�Z�?�6� 
>�z��z<�(�x]�Hu�����E��l`q���@�W]}<�~룘x�toBe?9N����+e�꣝/��C�K�昣C�B@W9���Թ-�럌��J���ۓ���L ��y5c˺'O����`AF1��m�)z������|u�X�;z�i�H�����*�ς!)����K�޽���;��)͈�(�L2v���J̍u�dsJ���쪰7��O�[��@T.���z���b��������r�sViG҅o�Jg�8���'ҹ+�fs�bC+=�dz��YVː���W�wF�^����ԡ�fc$N��ь�rT����y��]��" ���L2���!:h��B�S��e��?ͱ�舊eX�g�z��=��e	]���P���9��\�}jO��d<�%=���k/e4i�����	پ��|��?/so�uC�滰/V_�G�t01_�v�wĴ��i�d#=L���($v%5�G����6�mk�0��VD��V�`�Ģ�'�~$V��mu�*v����ߒfM?c4(_G���*��MQ��1|:G�/l�z�0�<�ڽ�.��z3$۳Yxı���x��W��tl6��` g7�#��S#�����������v��G�#-'�%�6;U�s,��W�{n�t5M1l���ኇ�U� <�ݻYw�*����L�2\��E� �����D����gL���zWl���0);�y�3��]��p���IŨ�F`��v��H��:�JH|t��%QBي:���}�;_l��:Fѓd���h���O(�3���t9\�V��,f�)�7]���ȓ�	�����!�	�m��\����y�������y@&a\vP�q+ct�B㬊�{2�8����ۧ��t$��sv�R{gK<�5x��8�C�Tt�j&��>�xzҐ7�P�
Nؾ�b�]|��1�{���z=����n<ԗc��`CY���N��]��9�����x��G�� n��4=r��!�Oznh���Y��2q�\�U�p��m��� ��=������T���'�gH�A�r3I4f�� �"P���C�>�>�~�A�#�	������3q����t~���?�ԯ��S��b%^�a���^�A�498�+m��tβL�/���,�4g.����Mv��f�	�I���q�-@�+��q��gF�����XIgl�dG;�ժ��j�EG��]}���H}>�Q�O�����M��rI�ik�`�f���r�G�|��$���}c�M��]�V\?a�[��ٹ.��ʺ� z��S�^7�b�~2��0/!�~1����sC���������|��,fS�	�p�����`��O��`2վ%����p����,�f8�0<z�fR�/]�k �o�5�~�	�T:C��@�3�W�开0��5�Έ�Z�Qh���`�Ͷ�ۈ�M�ë�
a�uE0�����̰����N�F��}�g�%��p� T�W�*8$ ��s�����U�f?���8�d��!2�>����9O&��u����nr0��RP�r$�Z�H��Ũ���q��j��lnT���8���^�/|���luïkUK\n���c;�a�z+1�ڻZ�j���ZĬ ;�q�a��y���8t�!2�K4����p���������������Ꝝ�>���b�@&O~�~�@/���Q��ZJ(a���� ~�J�(��E�~�sY]B+�ɏ��x_ݨ���%!=�I���g������h����>�,jɴ�� ��r?Ѝ�7rk�+�PQ�v�ep^��d�R�*w���?�G�C�]Gu�|4��}�����W���K@L��|6�A�P��L��C��&�4OOy���6�x�J_�D�8.T{�8����+� ��F����-�̟��[�/���c��
&ؐv��".��f���==/�m��P��L�
�oSHj#�M��2nE2��Y*	3~��͏<8L��`��?蟛��)���و�%ÞP��> H�Ҍ�*f���/�j����"_��Gm�w�H9e\SwT�T,�8��*�޳0��sZ#�m	=��V��	��K�\g��{}Kޢ�p�ٔ��%���6A��%R[�H�s+��]>�k�-�/)�T���ɚ�V�H��+Ĭ��m�Y�1���!/%���>����pc�%���/�=��6<���ٍG��T�=@�뎤�1Q.�
��3ǕN2��m,�X�c��#
�1�
��/��ޅa}�Yr�TGݖ����ُ���a�9�J����Q;��?�$���x����p��5(�y(0/���E�<7��ߟ��׍��gf��.�ེ���gs�У�FX����J�SЊ[l�s��t�1�����X������P�절�����3��Mz{��}�< `��`
y&R�J�H�_,�>���u����9��9���[g���n�R<�Bl�[��$1�SWt�%Ȁ"��'+��&�Lz�,�{[�-�U��PP�v�ـs�Yx� L��u;���Ƙ�6-�wR;e��s������5��c�w��ޗv�0�Ƽ��PAp��tC1b�޿��A�  8/w��_ZNu��#�B��"30�t
PJw�h� T�W �6�S`R�t#;:�h:䥎)��{����2�m���0��,R8.�|a�P,l#Y!����*��3��@�ɥnj2��������6!Z�$������^Adߋ����7��k��p��=W.��
�Ɯ�ڊ;��"qLz4���X"ע�~���j����@x�x�ͯ���㗁�2m��<(�Swö��,����uO��SIC���7�Qc<�,A?�n�-���_76���B9��&44^�s�J5y�����T;�S7�n?�J�@W�ΈrB>-�&�?�����D:�d�[�c;I���2��2y�E���y�U]x4
�P@B�1�5S�>�4Ƚ�i�Z�|U��p�[:�3k������H�u@+�NK��j/�
�@Ŷ$�̊���a5h�6��Db���v5&�r����0fw�i��5��g<ڼ�G�Ģ��#;�Ҵ��ʕ�3��ܓ�%�2Ԏ��6_��Cer�����rR��"��C]L`��ZP�X��K~n{>jh����r��N�D]Ȇ"�w��s���-&H�wO���c��a˿� ����ּ���;m�K��e�!q��˵QPX�ǒ%?4Z���c&�0��Fc����Ph�{Uӓ�j#2]j��f0+LP]*��s�(�{G`�� ُ��9��DА>�	e�ͻ�Abꐗ{�͉���+�5ā�z��!��mt���(g��w� �X[s?�N<͉P���{V8[�[T�<�(�{��Օc�!�v��B��:|�L.>\�c���6l��Fx1��Țр���k�7�a�|���c��1,�PD��w*�`xR�<���KV�1�3��2��|*	�O� ����h�L�@�w��@�I9���t� '���0�D�0d���������u%=�3ߢ�PH���W�4j܄���W������T��V*���n;Xvg���Pޫc,�ؐ��,V R v��A23�,��s�:�pzAz'�����SVi<?��������I"�n�+����{h=�?gԧzW�2/zQ��曠�I��ߌ�ýȗ��e	Ű��"�C*3�k �tc�yP���?Tb�������Y됂<��o���>5}����UtxH4��_t��멗t�&�od�3	!\�@r���V��N�0��m��i��w��b�á�z��ۗ�.
x��K�ă��#_Aof���u�p`���J�%�R�>K�����فƏ�B�������&����i��9d��{��nԔ;4'��1L�b4A9�������cO�)2�6/�����vfy�{`ώ��KB@�55�HZv��maҀ��d��^�h�l[�д�]�Ac���`% efj�l;0��Dǜ��ձ����Z��+p��P��n�J�ñɚW^�g �<�ڟ�pP�C �-���n��Ea�i���J��h*w}�v�	t�@@r�~k ���/'����j�kۯ%)DٗkG�9��gb���-]EW4$]H���*���Į�w.M���F�x�S��M%9���F�fx���w���).�6�Tz
��z�UI?an0e�M���.B,"	ڐ#ǴA���RmƴU��Pu5\�˶��v�D: q'�V��g ~�RUn�?1�&�Ζ��m��+@d��t� m�Z|�=��]r�G���
y�z]�`�؁��?Ų�u�s�*�EFL�O[��3�p�i v�E�s�T��$9���Ċ�L����%����&��n��ʟ��N0�W���W��F�6�C�t*yF&��z6�!P�A�^��"u�nËfή���_7�&��������e-���U�����V�z]y
ajC�t��Q�_췜�Nm�p÷!�(��*d����IKI�0Sw���B]8�s �F�)�I��9��n�*��<���B�|?�<E�ܼ��<n�}��{���2	fe�ĺ�X�>_�މ��*F>z�#:��do/�G!�%]t.ԜXP$8���6@F�#V�A�t��O��H=!�f��C~G��P��L���Q��i��.Fe�(��M�ZXn�ӓ�D�ع ��3b��w���
��pp50�~A���Ť����UF������u�s@�Ts]8�@Qh���"&��T�ܒ�R�?���{m'���qr�fl�^b���Aʱ��Tˀ��$�5:>���Ο���j��ݺ�Ip쬄��ESm:�N*�gi�}r`GP���S�rd���Lx�['��ט����քw�TҘ�f�cGq�+̡<����������{؇����Ҫo�H����v�][T�$�I�,�Ž,C��<��`��S�=?D��R��r�Ƃ�H}�ѝ�� �ڸ���O�%�J�L�Q��=���*@	�0���n��kF�	���a���n��H�U|Dg�k�4$�9��E�3gq�J�X���xP�@��Aý���4]0�����a���O�2�������]c��TB�UH{�]��Y����+;n�rW��5��0�N�W�%d���u�qKQLb�J�L�J
M��&�~'�P�g����q&9#��{���Ur�|��u�L��.G �ٸ�p8�3�`>���c�ٔ���LǕ��yJXٷʪW7|��L��`P���d�=�k�����'OC�ͺ#��� ��rC*2�L�Dx��K#�d��2��]v��U��jD�-�Sn��<j�5Xˮ��=�L�Y�ui�Xt���6���eҦ�t�49"Fs}u�����b�DV	�;�Y�il��
&��v��������M��������d�tWbYn���� ��v�>[Ϧ�~� K��BQ&��kl�Ϗ!�1���ܬ�D/�I�l��0\���o"�+�9) 6��L;�*�aW�h�h��E��/Le����5,|^ؘ�&o�|��3D�NhI �Ȩ�Y��Y
Z�����q��hkSM���� I���bӊb>�k$!�rln.&zx�{��/�U�mQ������Ĵk��8S�y¦�%�!�A�['��&گ�^h^}�!h��lN�A����]����8G	2m�v��e�NQGUT��$8'�Ǐ����Рf�mI6��|X�C�M>���c]:��D�8��,�/�_��g'�I�DGi�H��~��:=��;nw'E�E%��j���!�4w�d���x��^ͅ�{0k�,#�V]U��\���^��`f��|H[8=V]�X�M@��\�1�GNA���f�T`�^���t��ʯ��ԤDų����?r��*�� ����X���w��Vc���5�x^�n��,�q�zXm�OEMLci>�z�s�!���!o�pY�G���K�0����<�5w\㪢����	��o��(�8!��)Fn�%l��{T�[&�d��%��Lc˨+�K��*�=VT�� ��h�$/��Z�X��p�4���)Ǉ�����7e��o#j�zE`-���xlt�U ] Dܹ�4Y�G��^��n�C�Ui�'G1&��	�D[�%��o�T�=U �MV/톢��Rؕe��3jitH��b�M�("}�e��Tޝ7�i�2�A;��a�`�9���8f�m[�K�dΫ>����2��l��WZ��;���i
PL�"$��i�܊�A��L"�r8�/l�ϽLK|�b9�qؿץ���.9��^#�s ~ES$��Ԭ�����w��W�g�qU�tv�rk��0%���K����&[:�4̅�mx$Ś�r�O=�{�{s��H�M�-��2[o���aǽh(��4#���M�f��Rj�Y�Z����I) �{��*�]��Q?w��b�-��f&�O���Zk��?�J�R�c�qb|�ˌL1l�ѐ-9U��M�8�n�*�=4���D��ǆ����A�Cz��[_��+s<����]o���f��.��M-���mZ��݀6�~�i&	�?�� �B(u6��#C���$��;�ro2�ּ1ON.w3�#4�������x�8GB��i�ܜ�ym���ۦH�2���I��)2X�mq�!�~BM�/�n\�d[>��{d��a�u����8$4e+�ѓX� ������*�U[��~8�˶�{8Ǎ�6�QL,�a#�2�ȡ�TG�ع�ˊ>O)����P��WI�a��A^ZJHj���\\��@�Φ,���@��~!�K1�b�^/���W*��%N��7��'lBC~��}omw��~�q>���"`M�F����XR��q�	���
5d��e�+�K���s�Z������!Bkyi_8
U�����)���H��c�$����U�D�g �H<�Š*�i*p]�I����V$]��ɬ�Q���J����
��$z����>:��G��41�I��|[��A@��1܌k-!%�=3��MG�`N&��HFE�!��X9�[1��c]el������H��7�#��7б�����2�_�%?w���� 삩=ޭP���.��-���%��$�R�}HI��(�(gY����(��y�{ru��]D�-ɢd%��O"�2��gAC��n��)R+�lA/j)"z3J���z	D��u��O� �'����d!�0{rن���d�}W������ɿ��#�PND�l���)^b��E���ї�|;�������M���i+fyQ1�x���8�etƟ��H��?���<�&Ɗ�����d��e]>C�d>���&��S\!)�����k8�����R؞�Ÿ� 
�кE����%�y>/˔vWG��4p �;}�%,��_o�H��j��189Ǚ��-%^6��n��e�6I�U5�D����}+�$K����]��lx�����s�ݔ����� ai׫�I�?���)UK'��/0�q�`����Q�iz�u�J���6�#���������S�J
�;�:���0T�7t�����^��s\�j�*�� ���kHm�3�~��]����(��OԺKL�������q$T}*z����{�>h���>���ߴ���v��@�M��L���+Ts;=Dd��cE)�R��Ω����^��`��k�;�����a_%E]�'�䷽_��K���qy�h�%���n���O� ̞����-6�lt��_o�����%B_�%��9,�B�;
��p���B�6�)	3A��Qs=���ڝa� �E{l�+���߃��Y.�Ԗ���$�n����bi*���]ґ3�(V\�H\��H/�1UBb�@e
���#צ~�>��z�霡B��-�r�;��F�t���R���dˀ�}�l�ld���&�76K��Ds,"﵀�
N�����Sl��KX5W�E9A�[2���r�u�� 1�ڄ��-�3ua,�J�(^���jK�� �"���8br4_����M/�q+;n��nt~jP��� �&���H�A���4-{ ���7u����Q�E�m��%�ޤ�om���U�G�����^�tO����1Z���M��D̜�����Q���T�7\Zۉr��#[^�F�"t,磊�H`<%/5,k=�:���T��X��ӫ����ݾ�"���*wdAX����̶�@�H//DlY�	c�U�K-�z5炳�3��'��(���e\ ��b��{�r�1�y �S��x�;�7�nƔ�k-%~��֒T18���I�s�ܭ�`���1�����s3�-!>_���bt�� /��W���ʏ]ϐ"w�����bV"�.�����!���y�o�B�*&�`D�CV�W7��G�'ח�1ְ�T}uq �y��Z������~�<���"w����NH �H��'-z�A�-��p�)�Q����]�.��.:'\	tsV3t�zDO,��{��bpd�W�>�܌�fBsn,*^��X����|����L�fw�@���G�L�p�>��y�j1CBp��(
`8f�H�Iq\}�!쒊�Tr��7��fG�ߞ�X��j��MN}�{mI���ۚ�O�/B$����.б��Z��Y(� ���f^^	z�!�fP����6͖�W�����>��/�����퀁b@�0��=H�0��a!%�dS֍3��,5ktV[@F�����)��WM��Lz7\�-�+��ˋ��J)�i':�.\ڽ��Z����:`͂�P�?��\a.�&6�$	O�e�Ǣ� �]�kz`}x��I���@)PC��X.�,>_o�F�ה�;	�y��w���}/�#�M�P�S���7� G�L���\��% �s5M���7�,da /)�j���ȟ�-�/�u"$��}�Դ�#~?`o��d|b�_�@�Hy��R�>������ƫ�`o0����C�׶��]���ExfG��T��>@G��'���髡��%dB�ϱ	��j�ZF�&���9��R�Xr�� �7bq�3�A���|gQ��֪L�?� �G�$�{�� ���P�jDn8�	\��㴁O���������ًX!lmy��Q��Hs<������n#S3����G5��w:q}�5��J�:�_�C#�m�������]RM�*z��أoGA�[�k����C����~�%�������6:�K�C�W�І\��^5�bnoP��ǫ���:5�rߙ���D��w{�Y��.�)9(�����������2��>��~��7ˀ�'���U���ZX��r,����(�N�e�|S@�9(n�jB��3�o���;V� ��r�Mn��Ӟ��^k��%����;L@�����P�Op����*39 � J+�"I�|�,0����.\��E"�-C�lגi����x��U�� ~H8)1����"�-��0q�{	~h��]I�-��������X(���c��bD�)��G�p?�v&���sX}JCYv�BB��lg��X<eCㄍo#{��/�O��DS���T!ˣ��7F�ئ�S��������Fү~���� �Uזۊ��]@�@)��-���|s�s8{4+Q�ܸt����e�w���am*��.�F=�L9\�����?˚��`	��yU:�u����l�����w��\~{�ťG+����/]om� �����b�M�&ec��9;��� ��`E-2	Vj��)� D�[�t���0VX�%?`|�������f�.�$$3�R�=c5�6,��l�(f�ɨ���//*Dd/���5��R/���Y����뭲!��	�m.��]'�.ut x�jd����v������|U�U`pKY�yQ�~\7�>��~ƨZ�Q��S���	4���xL�݅�r��(��4�.h�P��/@�ǂ��I���Ғ��lܭ����%�τ�4>�Ȍ��t��`X�D�0 +,�כ�cl}�)�v�^��Hrmj��~�S�����Z�ӎ��0�hqw n o߀XA�"�x��FM]��,΍��k/����$$�U���3L���?cڸ����wj�&��)J� �)�V�'��/f�$����B��-�v�R��L�i�'�1vF����b���H'�V/�|6�-��z� ��ٳ�l�=SE׷Ģ���AMo��^#�����K��&�ַ���ǋ�
ƞh��q\Xqg�ĔLy:��X���J{�
�d�n)r��]+�B,��e"��7��p휳й�b�
���L饱�:�V蟉�W ���i?f /�D���X����h�9������)a�&=ʇ�}|OM��𛏺jl�s
�dy'-���t����xɀ'FJeˎ��3�Q��{�1Z
����*�ϗ� �5��.���"^����v1�����ˍt��m*��&�Z�`ʫ8�M�r����f(?��S�8A%D�<�Rfia����^�nhFz�pjԤ��p�A�f)����Lv��K��$83ʬE��n�J�C��H�K�x۞P��9����s[�X�uf�;n[J.���C� ֕�������x�<@��|�@l��c���fB�Y!�c�c�
�q\J���p����;� ��n��lBS��޲�k�����BBy7h/��$�d�B�_W�����A� ��S{��HO�5���b6y��~1�� �܆�ڊ�}��ɰ*L
�4Z�� �E�ٕ^�n)�2h²�Ƕ������[u���j���Q#r\�и���#"fI�sQ_-�&EU������d���E�p�0�Nn�/ؐ��P!����2���>.�Sȓ#����Y}
Y�ÑSd'
3��W�ţ��;V��&3�I-x��L��6����������FF>Z�Gi��E�1���,���M�G���r����'��#�PPi&��c�Cq�\�8���Ȑ!��:������A�A�п�V�&�n��e\��ߩ|Ï�l�V�Ymj^�`c� J��d�-�=��kez��,�%l�!@O�uo�����nK���2�(�?��%G��
�-��g���h�	y�Lk텕+Ӻܗ^$�a'�K�@��綳�{o-C�р0oŃ��u�n����F��o�6�Q�P�?���Y�I�<�Z�qe�q3��{5�"!�s��!���8�4�|Ru��9�6���Iv"��r2m ����8!$� �}����~!N�x���ޯ)|���#�l�	=�}];�մ�t���@�Rٚ��V�S�{��h%�!����V����y�}��8̟;v ��+7qk��"�H�x3��1�{i6�掿�g'�-V*��7�,`�㜔����Mk�Y�	2�Ze�/�g*�T͐PԫcD���O��m��������9���Zak��ppm��ю���������έI�U��]K�L�[A���k�j#[������q(�<0%c�͚����@o�Xq͡f��`���a�(���_S-E�-�z��q���0�I"�c��&R2@�p<@�iN�qߨ��xhCh�1x�k���n?44�2O�	D^~��[:�E��:��R1�taC�@��ta��RN�-����p��ԕ����a|����v�D����e���:Fx��IB�%�D z(�%��4�~�[J�тo_��;����a���R#���q2�:qU�+�U1�e��rȑ F\!q��Pp�Q��.��\���B�T�������Y6N9���O�A%:�=�e����$gwt�>��̃%��Smr|
Y��<�
����g��o 
���
�E��oZ������ֲ�++��u�� L����9���L5 �2�y�c@~�'~o��~m�E���n��dNX2���`=��=���*�����r԰�����/�_�eCM��M���Ѥ|Q~X�㞕�D���˃Y�º�,U֕%��I
�6e9]���:��&�Գ�h�kO7��=,B�&Զ��d��t5�p=����#�2�'ePg�G$�a�T�'kq>m7)��D(��Įǂ����cw.�%eH��b���Mech��WͿnu��NTxt�B�*�8�`��������v�܈�l=:�Е�)i^�烺��p3�;_@e�Eb�p�����r��ii����Л�i��zQ�h5X�z.�0>O�ю\�4�"�U���?����;�{B������� Z��0�a���Vs��L}0�?�e�q�5|�vZ�k1Y.8��W��8���	��\E,��B��0D�{�&�S��OtWo�;�ޛ�F����r-� ��'J��%G�@�nj��=qG,�FSJ���|��7�. [�z����X�٩l��*h�&��c�W0_�ڬZ�LJb��N�����,"9��8_����(
�*��~�_,� �c��Jp�+L(!�\�!#�i4�'Iω����wHv�`�͌�� gU[9����,���B���_	���i�s������,�Ū40��0^�F�+K��^֭�$wt?��yZ��B�lNU�]��fU�26o��=6���k,mfJ�zDf�$�=���h�p�h@�u#��o�)��뇹�8=ؖ:�L���q��Rg�OWz����TeI��-?���\�e:��A�}Z5¢^�T�s�fdQx��:9�UTd��#/дyktn�mN_�*���$�"�<�(۸��2֦�u�~��H=�����3�b��QP���r�I�0����a �z#G�0� G��r�W>��� �J���r��b5p�~���н`�l�,� �i�r�8*��>!@�oX�6j�L��Q�5�Ј��
�="a-��N���ZI�I�5�G��rޓ����&ʱq��,A�-	�Hs��Y(�?� ��^N���֫��Π�e�eQ�e���%��n0�YX��*���s��J�;u�,U��H���qC��
b�<�):�Ѡ���v��Xl�^1$~'�9p(7���>qъlb]�>Ս����qnY��"��*����5,+� ��Ϛ�HT�n�1)yG�wj��y2�����'d�!�q6��6��y���Ha�"̹&�������d�E#���Y���.{�x�T���S���5hx�� gϳd�x|?�b��Pi	�B�S}x:�KJ؊w���eOi?�t��x����x��6�Fo�v�j�#��击}t�Z�F�X�����C�n0�	�x�HRd�zY@�WSa�ț6���HԦ֎읊5��b�T��������tLL��q����-&��6�u���()���,,�f�Q�ߵ��S���������B��-�E��V��>`��8O�iͧǠ$nP����²�I��#r(</Ge�q��@�NǗ&����K���4�ĳ}XJ#��p�A�d�NY�ٮ�\�ek6T��ԌrV�W�qA�^/SI�za�z��%g�nP�h
�5��D�Rx�7&V�{��"��U�车�h6ǪG���V;8q����j, ]���f*Y��xz�a_`�>�����Ѧf�w6I��#̫!;N�;��PzT!��٦871�7����jt�S]��f����8�����^��X1S��i1��OG9��!A3N�R�����1�x�r����#�a4+�sGI��?2t��6� ���w
��ң����c��ɏQ���]�Yı��'� �m�9�R�8�X�����L��cƯ�[�0M����Ni6����r-���/��7G��Q�R�G�Ɯ�L[��G���V����\�E
N���1`2�D��.Y�y
�L�p�|�I�Xð�c*|1�dV�<��n	�����C�7y���j�9xOq�s�[hp�q��{X�`V���d�e+�TxS!Ht��ߊ8�|�Y���(�ס��p�-�cwi;�8̀����Z�dC�et�r���T8�p?����R#|�v(#=�"�ӳ�%��0��+8239J�s�.�-qǓL�[�D�����ٌ��?�f�WA{;�K��I|zd����7m�M�e�t�5��5�Ez�K:OQƇC)����5����d�����,y��~~�E���V��V�AgN����o�<E�L� ��Տ�����;�h�����~s'�� Gmv�A�D��Ə�>�L=���&�����:���:��؊�ܕ}|ŮD�}[U7
�1�r�_߆J�}o���� x�qP�m��e�F�1���Û�Sك�o�dt4����6zT���B�f�}X��@��H�N!���ckS�p����G�@��!WQ�fj��|�����G-���#��|���oP'��BX��ju4q?�٫8���U�*B���ї�|�Aq*)��62c����|���ge�@1��J\ �,�	���I6��>�Ә��>'e��?ޅA𰞍T`��3=?�(_�J�qNT��l)p���Q�[!�f���j2�6^���!�QU0"����U=EУ!��z�f�v aM/�x�(���Ͱ���gH��箚m򩡔 %�m�8AnΜ��D�V�e�>�X�(ϒZ��D�R�c�'j��߆m�������tj��D��Y�T C*�����"�.t����]��a��d��w���-e�Rɗ*+s�Z���w#����˚���p��I,'c�;��{#s��V8���cʤC�C�cJ�B�<}���gM�;�&ܳ{6�yM�pr�^f%��&��=�(kos���W�_�L�RWj~@�ɫ���5?>4�p�MgQ2GU�9���Ϲ�^��UO����*9ı��a��L���a.>��8CbVN����\�u�8���!�6��rIb�?���e�c�|ј�,��S<~�Ce��s`�0��>')��^t��$� f�����0�`p^�콈�a�Lȇ�[~)
��^ڡ��ix�B�����m�B�.��N�}+�#��}����K�~[��A^c�n�0g��v��L���5��a͒�o@�I�@�#������m����J��L���!�^ˆ�(F0�Wz��g�J�4��MϞ��A���+ʓ��"�A%��ȱs�4 ���I��:s�$p�:jc��r��'�.�sA7!��� ���z<K�\��RD@]�����	�H���G�1���	�v�u�\�|�:��>�'&3KU���;��Ct��~�4�8:��L��L�Fd����&���~���NW"k��58�H̘�;7*5hh�BH~�(���S;�x�ڋ�$Ej_���2P�)�}�-�qꚀ�2^���$v�.��N��G:������@�${�t��[�� s�0��LM�1N�[v��m�*"�m���oB����@����d�3t�${��;�v���y��xU.��s*9���o���w/<H�sd�/���5w�J|A޴5Y���iz���
9�bA��i)sX˅�j H@gb��N]ǡ�e�* J�(jYt�h�㰃dw}���/>:���RI�n[���0*�=ۊV��-�f�/�]N�wh��-�1�7�me��!���:���3]0x��'�V�&���e2��(�;�0z:����.��h��ޡ�@9*˄i�b._]�'ܙ]Y�"Kh�Hll)V��r�P�W�P�Ř�Ҫ�{��h���T�/`�]V$R@z)��r�	��]���4"OȻ���L
�sʍ��7-,�����""Q�U�.���Ȯ� (Eo�3d����{�M�X���P��T�H�HPpI��Ԓ�%�qw��	/ȅjQ�7���YF&ֱ�H���MX�,����z��1}�g�h�-q���J�'��,���v��W���I@�� F�����d?���S��Q�	�~�]	��y(
���e�ؙ��q
bX�u��&����W�m�$b��V�Y"�34�.W��r�U*&�X�GWU?�5�e�S�D���ǖ��7b@9�ޜ�-����8��8:�t�|�4aWY��Q�
���G/]Dۜ�Kea/�� 9�Y�#v�� �6ό3��eM���쉿h���Ų��TZ,�#��b[�4r�d`��~����%.BK��P�'�>r������f�X���$P6�e��\p�t��qD�����x�\Qb�O�����±��%�ߞ��wy�_���V���$��Of�����7ƀ��%��H������&+f� �^`�st�X$p�C�}e��t"�-^S"+&���+��@�(���(G�]��h��n$8�:=���%�9p�q��n(]�+q�#�$��J��mh��J�c���Tf�E"?U.�bЫ��P���R�'�Q�&1,�梑�L�3b���l
>�'J�D�r���4�<3�9r���*ދ|2-���U�hM���`�`�&�$����p��h���=�9�Prq�,�88	�3E����� `��b��j�$�ޒr�E�����O��{���SDg��oU%��@Fu@�F
��I<M���q4F$+
������>�w7S0�5�,�N� IF+���D���,�>Nܐi�K)q����d��H�A�\?6Eg��1O
?�2#�g4W��]3�� ���X������IR������,!-oJ�95��ƍ��x��Kb3��g�X	Kk(�EAT�h��tu��˚��a��5ZPl�n� c'�[��܈ZXP79l��mb�KLA�/�����t��j2���^�GCh>� �ۺ�\k㞫�Y�q��"���n��yl�t���x�i�;��K�,����ݍ�O�?�D��t��&��&�M����@N���i�@�=0Ԗ;���g8���Z�hJU��N��cr�Wޭ����j�&:o���9�T��7Ho��j��.d������^���-����f#Yon��E%�<.k�M�S#� �Rl��:�u�<=*n�����C��J-<��)�G���CG����(
�[HX$�"԰Y���́u�%VL8whv��ߠ�=�w�.te�^����c�4� ��+0դ_W�'��ԞjaK�c�.��Ja���E��f,\_�����m�C9��Y0��|��2!�N�-���ߪh]���'�� �Z�PݧG�T<����F��z��FOo��IB�Tgn�N&�L�\�CiͰ��M��Ng38\�&ȏ��T-K�'�<�s�t�ݢ�m�րw����RS}�c߱3�����T!'Q�v	��#=�I��3�|�au^�\�XΨܴc˕������ō�#���ܰ�.�����l%�Y{��D�}�]nA
�l��4O�lLcޱ�~c(ۇ�<W�dD�^ۚ%��Ռ���˸w�W���c���&R��SD����UmCS�O�a�4���3#��W�A+�^-ŜAJ�f(ȳ���U)C���c�-�m
�4��&yHAى3�+{m�ƶc���s�O��|Ҧ3������ϐ�;y����LSL��lԹ�}��a���p0@�ј��?xء�'F$�S�m��4��L.Z��X��X`%9{ë/���GPYR�ao3]rj������d~^��b������NV>|F���۸��� �(�D���x��T�,o�� ��9��H���q�Oz1��1N��3��R��ӽ�a�wZ@�Mސ"�� �R��I!8.sS�y���s�P��"��%�*�/8��֑�<� ��*��*Zx�}���>��#���i�$����X% *`�Ɣ��WqG�ge���x�y��?ji�p0���^��Kg�(�����s��&Vo���K:�(��V�&��9�:;��]�J�!f^n��iy��8e�sW�@n�G�b݁���v�g��f�D���j�ߗ��J�}�����=^\��A{o�(�qd��γ�y�&m�\���;�{&D3��7=���u���<���KR{ܮ��˲�8w�e vnPȞ� �|�E>9l��f��JИM��ĊOv�4i&���T�,W4�D{��S %0��'g^`&�ؽ����F�1��'i���F��(��Ց_1`�D���f�v���ܱހ�5AR!�L��1�܌��.�N�@vz�y��(&`��K��E%�3�O�|�������g�Lȳ#BD6�4��wxj�4�d�A'^�J���*I�-t��䁲1~iK;�Z-f�.=���""c)��a�y4^)�Mt���!>���gą�!����=9^�{���j���(T�]+����:��eO�;GP�A���ڶT��+--�i��0�x�m-:��F�4)	��8)�Q�1�n��'\���g6�h��a��%T:X���{\�P�צ�t��m�ʁO�&�A�c)L�b?D�$T=�=·�N���͘���*>~��:5 ���X�%������{��P���f��_9YzR!�� ̚~zI�����A��¡.S����w�"]�,V�)곗�Y��ptS�˙�f�ZM�j��5��<�9��t
�f�x[��X{����7�����v[x�Ѱf��l�qVC$Z� Bp���B�A�23��'^e��4�� ʿK�g�:7�dv@�Z��D�j�A�g̎Tl���[X~\���$�����bK�ԭ���{��|H��K� �SO׆�)���	*b|��һ���Z3ua���1�W��A�t�[����W� {�%�P���y��c,��q�2���l�f���#,"�n;D�类�U������d�#�_E�&���۝^�%$�$��v�2�`�2���F�H�S������ډ��./|�Ɖ�\���}�o��E��K}͉�A6X"�~$z,4y(��zd�.���
[;!�$L��F��������c�B�ش�ւ븮w�ʦ#߱ʧ5�~�`��p0��YC1�1ĭ���I�����(5�Y�<��T'p�����n�^�p��8����R7����!�b8�ē���S��:>➔��X�l�z	ˑC���������!s��(���\��t��MNH���&"� �l��ɍ�໯!��]���%5:]_���]kܑ$�&즗����aK�����)@I)�-�D��Ot�Њ+5R�ѵ!0#(n$���� nFD(�}0���8R`���[-�~�Bw	�d�����{�nZ��ڢI�	?�4��Lӝ�nff��E����+�����֌�ԥ���(۹�@�k��'=q������7�j���h���_���O�4�����0���9*��t?��?5�m5�$i۟"����K�z�2������&?`.��~rE4�01X��3;��Q�1��ڣG)\��&��F����H˥Qw�X�2m?I�!�|�� ���G��y���)�ۚ`���I!��; ls�E�X�c��k�JW]���n/A��`��N �u�d�d��@s� ��&L�������������2�t�3�>�Սh̔��S��� 	l��^HICu���K���ɝߥ�fֿJ��ң�m<�i������9�픪5}��G-�B�s��Ȭ$P�U�S o�G��@�އ�Ld��U�y�ѭ��A��͘J��7
ގ��R�����x�4R:�M�2����	��������u."f3�= ae���O�	�����押�|&7��Ze�2B����7k`���B��R��h����ه��;DW�	[�����a��࠲d;��Zܞ�.�K�uoƑ�q,j�
��C���'��2��i�IȎ��wz�ُ��S�؜U�G��k�R�/Q����%S�������`�&��`@�>��oKw������Ȭ��(��!<�/ޜ2V�Q�eP�۠��4�)
��N�W���Uc��(���r��tȫ���E��{-��ϙ����Ϯ1=I�M�ĵ�+�����_:���$uF����X�q��e+ɳƈHkk��]-��S�m�6���֥�9�ֿ����L����;'�bn�K�c/O(�˝�*��}�mZ�ğ��'����j0���,ž�޿��ԆL����ܛǐmXx�=�r/��N��A#�ϴ������8"�hN
�'�����K3���e�Li���믭'Q?�-$��oE�7�q?�LK9�~�#�c����!˛m/���^������D����O�M@��n����
f��y���hF[]��=f\Ó�1>����P���.�A=B�@^�E�>"�)�l���_P��@p0���0س�cr�D��a����1�ޱF��y��`���)��RA�i�Qb�5S+������*��@�:W8�~�ذ<K%짞�hb��D(cJ%�֦�Ae��	��ϛ;3k�[�~�q,�,?z���}�n:E�j]�Z\,�j/V/5�Ɔe�fC�j?f�q⤲�����ʚz�[+J��-v�L��\둻���l&�d�I�4���U�X6+c��0�a�������W%�n�i��QW-�x�D���}��T�v��o�M��*�͖sJ�ei�iYƯ�)�X�7ߙS��F��X��V����+ѫ7��&BӍг�Q;��8�u�x-ȓR���?\3�g�h�]|�I��x�8�uvi@{�9;��h�O��)9(M&� �ѡ
�K��-�tه���\����#KP��v�:?�TRF�@�5Զ 8�y	�� ���W�y���)t%��G"d�H�Z�������O!����gl-����X�����'��㓕��5
a	�W���t�ܭ��m�6�гcÒ˅�n��K�H*幽ְ�p鷦oN�+&�=�Ѡ`_�h)z0kl�.�H��8�����ޥE�V|2eO�Y�&�o�qJ�����%�n�50��y2��<űj�4�ib���v�)�>(f4�Q��m��<h��ᕭ�����X������]����H��6�B؁�ue_�Z`��]A4M.Z6��$6��lv�q��u��l��v���z��='�ڻk���:VI��rK�N��)�a��� �j ZwՁ@5龴�d݌q�&oº��9�}ቛMY�����Zq�Z+��,�<ۚ=/\!�t�}��-!��9�r�ALit\���S�m>�W��_tݶ�x>�/ƀ�	Y�JX�7kP$�T:[{}��m�I�Z����c�����z�L�Ai-���4'#�|5=�������˟��g�A^���7���	v �ɥ-���A''�;������<b#�*�i���<&���F?k��O=rj��i��"����0'�A[�f�L	J��N���[w�2� !SM��!j.}}5�*�֩k�ka�d�G�{*��5��B�(2h�'1���|��z~|(1%�W�amkQ�@�=�,��c���Ĥ��Ʒ�T��@��B�dp�I�o�yde�G��:��(�?DߗĖY+�#�Z�F+�0�p ����L?I'j.
����q�G5h4�F{M5��+ѕG^k�:xx��^r�{k������+��ϗg��0F�r�����·��`�[v4�!��ja(��A��S:���td��:D9ͩ�&/�j������ԛmP6OX	�'�8�
���z)zY3].�!a�ބ�&Sq�y�M3nF�o�nn�넸
��yhnsm���3�q8�X�', ������&ȭƑ�	8g�{���'���h�L��0o�t<.r��g�C3���!?�@��k�<7������	l"��˷� ��M�\�yX/�ZH�_����xC�� :󛱅m�l,=gq㎎$I2i�^殯<���i�t��<��#��3I�Sl��]s��w�%�M�/�I�,��hJ�����"��e�Ij��">��]��b۲�X�������G�b��'g�W��M��Az
����ф�c.�:�)����G�������hjBKa[�3o�%,b��wG���:/�CL;=��� ���n`���;FZ�����q���	H;Z�XUNI = 3�x�҃G���E��x+uB���ɦ�'GNh`�.�C��}����Q�	o���ź�f�����{C1���RK�MyI�y�S��.��vL�p�ʟh�;���q����
�@�p1% (���bD#C>�8��(�z�ߑ�?��G�D���T�.�%��Bu�Ƌ*�[�����
�c�(��J6��OK2��P��&'�����5��:����������]Y����5rD�-��uDd��H�V%ņ�s8f��*Q]��ɲp���D:�J)��Q�c����I���?T���pB����4}�	�O
�^b��}�+����;Y$����+��=�Vu�σ��횹��~P7�beu���d���6y��x�4�v�G��7���P��v	Rb
"��u�����q4�3�N\.K�m>jƅ��7_z�$L���(_��u�.��)汬�,���]8���ș�ۮ���Y��6Pc��x���|e]���6H��~�W�XE����Ď �Y�o����H����Q�5�"(��3OA-�M�#]aM��}(�Y;���/~�鞝BX%�n�K�\Bu]�g�V7��l^�� �fP���0l����M��.$�5�L�z�[�3E9�#���as�w;'���dD?Il�;s�ob^�"�y��(\� 4[�䖕�?^�[z����)��`X2�U��������P�}�meB<�"��s�iP�ߺ��]�[Z�Ȍ]�Ǡ�B�/�8�uu�_t�kL�4�n����֧8l�05���@��~%�i�?7�+��_��z�(���4�X��t�8�ܫ_�x�5=�D@�66D��WCZ�"�`�Q�'Ŗ��G��fI�+��6 f[m����Q��g�gI� Am܊G�"ͷx�W�:#���>̩CI�^�,c�0�aq
z�O����of�݆H.��.�&B�ۡ���mhs���h��^#�������-�h�Bhl��Q�zy�`6I�Ӟ�&˟�Ƹ�t�I�L/��;Y�ŰJS!��a�N8e�t��X��*0��Ư�[N!K���A�v��fP}�j嗞�S�1��F������^�mt)@O2��3�L����4���G7^���A�����kk�y�W T��u��9u���J)��H�7a�*����JC�1[��|m;���+�k�e�?��`�����D�Plȱv���'q'Ƶ����끷�v�gk3�I��%�P��J��o�l:�O�U��t?5�f.��� ����k�A�F}t2 ��H���z: ���'�z�Ō"�8�Z���0� _6w0=�6�8���TOy'���ϱ&<=U�S:�^%�=���ݝ〳����e�6�Y�ڐ�҆P�|+<��=���G��A,j�6=H)U�?bԊ�r���{63_�&����XՖF����
U���2N3D߷?~�Țl��|�B�~~y6��WJ)آյ�ݮ_�:;�=!�����=� � '?�<�o>��n���H}����w���H���s�?����wB�VI��Y��1<��oԜY �S�̜��DBU�ыHS��d������NA� ����O�&Lo�V���E�-Qt�6�͆2g�Z�R�A��u���7��B���cm:AU9�_��.i�1�V��?�2C_�5���:��ù|k�=ץց')��>)�R�b�� pUy���I-5���[���'�� ���V�<�ل�<5����� o儋�V��9��Fc�:�(@��+?�F}S��C�Kd�親�D��k���Fn��	.!��T�t�`�k�3C��Mxs���m8ǥ!*B���"�D+�ݬ���cEN���b���n :_q��c���i�[�i�g$/H�ﲸ`)��!m�͓R��G���a7�����ud�3c�,�"5�ݰx��"���g��im���Z�����������Çl��'��.��sNܩuE�>(�@� ��lG�aM<�m}��:Ӯ�-��~���A>�`���'U]�i$��3O)/�~�*mk����Ү���	L �D���>��(җ?gM�x�ɓ����G9�����r`��>R��~\Q�@�+�R	��рG��ܽ:B߅���!��{�O���Y��a�L0�P��
��P�Bz�5N^��a���ǽ���]��v��ܻ_c�X�];��-�G���3�W�|�oD	9_"� �2�4h�M^��%�b�cZ6U
�uzAt����a?z��E�业�������B�4��O��M��b��mrc�A�t��i@�w����o��h @ᭆ�G ]�o��J��� ���##^�X���hQ�3��R=D�N3���ζ�+���^�]�J@�V���vw����_lJݥ��Z�V��4��L�%�vᛀDe����"�8l!�|�����|�>�+��?���px��Ff1�j�uVML�G�奚�=��z{v_L�}x���4����yAZ7J� �� y8�zc2Jl�si�B��QT�)'x�'=\ў�[u���+]W8B��n��z5k����"��� ������������Q�D�p��y��1��}�Z���x��Ibq�����,��L�c��M�e��F�׊�%����N�iV����a���bw��!��Hf	�B`[׎���ޙ���yM�+��g�ՖmN��̺#���zbߙ�}���H;�o��HEYf(�[sU��$�X���hZX�o�OWq���m�vD�~�k�.�:�hg�r�)��M��O�2=̑�gPh�G���kކ��}�^8� E����	��T�-惆gahQ{^���NH �/\�e�PCz8�}l�2&d{l4����f�s�{QW�P��7�>����?Ÿ�!���-	7��R�X��l���b�#�
�b��,�x?Q� �8l�l5����3*�/�"� !l�뫩�����t�z��_�a���*C�6��R�W� Zf�+8���,�2��.���w���{l�1&QWŢ�7�#��7��kWсv� W>��E����Ix9S���ʛ�7��+ڊ������Q��B�s8��& uͱ���^mK�iXl�I�J*����m������Ao����+�6o����4����W����9(s��3�ܯe��G/�B�l�"�Ò`M��3�=���ɀ��!��Z��)�3S�={?S��.�
7��G-|5؞��Ҝ�B�P�A�M�:z��`��80��h	E�[�t�g�N$�(`��B!�:�V0��S�,7��la������*_�"`�4j�-�<x�����}3��1-\2��D�k|���EF���H�u5��������v����.sU�s��A��|^Z��=@�����r�o�s!1m���E���8�io�E���E��RPE��i!��R9*>&&�m��E��V��T��T��
���$>Y#�(א�G�(g���$y�&qKC`�PK�ބ�r��΄@��ɛ���A�B��Q�㗶�F�X�Ϭ��ߧ���)��nPR�<�P����iɆ4��V�20��Y�1.�L��X_�9��<�������]`0�˵aa녙E�����Q&xQGg���Ԣl�EJ>��ȅ�c�kC���O݊u5��H�l��0W�f�o%�J���R|�R7����^ܰ�"!�w�O�ad .�Ӱ��J�<�U�ۖ�_��U�c�A3�4�y���]<k�[���ΪC(���$�G�8d �,���`G��O��`Yω�I�↣���MH�d�k��m�X �����KH��ޢ�#��y.]�;�q����췍����olk@��vɎ�sDZ�h�Bq�J��-'��y8�ѥQ��Ӌ�o��d@BX+���[�[5�p�@����)��8��o�����w���0�����8�x��7�P?�n6���^�|\���m1��w��?���ᆴk��(Y���dې�M�Y6���5�=�k���BY.�U(Am�w�*�z��A�w�ώ���`�(���~��q����h��+IBcLZU7�=�1@��9{e&��3݋i�Q�oK����j����m��yx�3�+$�bת)v�(���*�nMk�'�-�5���w�����Sr�+^�����,���_���\�8��$�rX�&6��Kש1�*s�n����~S�`k6+��+�	����0���~H�.J�|pݕ� _]�����C�T�W�F
A{�����خ�l&x��F�N}☇G_@=�{��1R�~�K� :��^E�j~
�B6��U�E���-��K��)4
g�JF>�5j%��1��^���o��T�`	��fߔq񶬳5�|�I��`A�v��8{�ˑj��H)i3�00�6��O3nEtpU��#���;���Vk�9���(u�̔�T=�H��e�UÍ\>3�g���ۛ_�9u����+��+J��y5>8�+��6g�/+��
U�5s<C\)�]��*g��,ٌ��!�ӊ�^�S+�%�'D��D9���.��j��C0�n�ZYoA&>P���aF��"֞/�'��Wx���c]�.���`wEc�F4,Lx��ggr�O$��}�т��U*
����ȑ�Z�bQ��(m&���o���#.n�������at�{��]���BR��7)�Z�K9��X<Y�M�� �wQ�(�ٴ�d;N�{��g�>�=�휯��$ �C���Am7�
壶����I��u{��G�tM��u8�։`Ч{m�\��M�1ґNc����x86������N�<�2$�Yێ>��v����yW��9��5�E��,��io^*F�8c�h��-c9�����!2��b��������i[ `>����jV;�R�T9ȥ���\P�W��k�B��z�e��^t?�]��E��1B�����ЋA���v���ɻ�"{�����
|HZ��Ѽ�a+D�onLv���pT����!A����Dk�h~�fKטLG��-6xy7� W�����n�ٞK��
S%��}N��}c�"�&�_��ȭ��@K<�]�F��6��1k6|�S�MG�%�
������Y��/����'�@۔��	r*�'�E�W잊�����Pmz�]Aj�&Z/d�v�$�>�u���i��b<��괝�)Ű#$��N��.OP�rrG��t!u�5M��lt5��rB���7yW��L��Uy���{�DͶ�j�Xiѓ��rJ6�%�~v|��2$"skS��`1s��GQ��d��I}�0J�ݢB9�� ��&�^��p-��핽 w�.��D��pq��?R�c/��R�����U3�-ڝB�8Z$&e�l�9w�Ma��	ǤU�4�Yq�,t�+Iݭ�!�^J$�X��"�𥾞M����YO�V�2����e�����4��IO]�,G⸜��#�o�v{)%R�'����^�kd[�ρ_ҡ9-�lW/�g��芼%Je�$�˹ʍu�6i��s�N5\�� �ú��I|�i6v�AKÁ�͒��Jx��z/YN�Y!^8gG�ž;~�lR�p��j���Qi�!^�/f��؎>��,��^���z�cK�7-���SD^�hc����R�Z�,gN-���c������ol��FHL� �413�R������2_�,��:-%d�]�%��U�J��6��	5b;�� �����Ω?���&x�g���&�����"Oj��s�]r]��\�C����).Ȳ^�h{kcNdb���?��s7�l<�j�eJom�m��$c=:���r�i�'�>�+%�=�Lw뎨�X)�5թG��,������B�]�쨇�c�I	c�Թ����(Ҏ`&͟�R2��{W}�Tu|B���O�G���Yא\[�������� i���ɾ\@��4�X��"-���>m
���m�؃P���/O\��6A.�c�g�e�t�:)�d�2M��
M��hČTy�.��A��l��ӂ��bJ� �e+:T��E��^�E֙:�^��777����~T���{L��R�nJt��j_�{�T��B-��JJ��&�L�1Z6;�k�A�Y��y���ɧ����C�\�s�b	.��Q^Rk/y��T�!zK�!y�]���YB�,���߆�xD��o��pr]��|g�����i�J&N-,J{���r�tUcgO���l�3��`]�)"��D-m���9�uU��p{9=�<mڿfެ�1�z'�����l�
�f@ȥ�� M����rZ�����ҝ/����v��,���͸Ґq��Y���b���u+�Jx�slJ��N��4ٸ5�i�m,,���/ш:$�ڽ�gY�3=���Vx�	n�˼3k���W��4�"��Ozy�9��M3�������U%��h]����c���5ӳ�]����*�o�{��Z6 >�p˓������Y���ᢧ��@/Sv��௷H�
w~v�GN.�D!�9��>�ȧ��z�c+�9�{��F����PDw5�.i��+�On϶桬c��b� ;�����=,E�$�7�z�*�R��Mo�Sb��w���b\��r��:)%P)�X��(X���?MrJ��6_�=����3r��%skLNA��^T��k-c�	Óv,�(J@���Ӫ8��c�MI;^��&Q�9�����2��X�n�"d��yI���Q1oL&i*M��ٰO�Rq�m>T�I5?����g�����?=�s}|yz�j��tcROA�����/ ��
������g�U�U�X��*Excơfi���;����%iHU�.)�/t������eз��d�RV;��^���k�Z,븂�u��hB�p��c�)6 'Ny��=�#"�g)�p��;�K�ɐ�V$���8�n����V�Z���5�m�I����ë��kF:ע����G�-�ȩ�n�?�2
��������]�A׊�����Q�ԫ�?%1д-�?άW�4ħb�s&�u��T����~�
��OS�����o`�E�!�c
5�ie�a�~���.R������מ����0ܾ"3��z��	��̨�U�č���F�)�4��N�W�5�̀C��#����8*�pc"W�Q-�k�e���Tӯ�qT�XBO�C5��`F����3��K�rS�$#7Er����D�xfI�y�T9�E\�2�"A#�G�*����崁����mfV4�6��w���~Cl�� ^��l��|K�#F��,����sn��x�V�ݰ��3h��������⫆#��gy2קx+ݝ�*�!s��OD@����q�5$�o��B:6�	pIh�l�>?fy�Q(��܈
EHK=��t���[�����e*-�`�XE��u-�bw=L��0�D{?�E��(����6M����~a|�7�^M�j$���=�o)h��N�{kQυ[70�@1��v�B�5����$*_�R�UCj3E�r\�&M��c�6oL=���^z�1�&x棰X�P��F�p�W5az�%x,ϯ��� �ܸ�H�q����t{��m�O�&���c�]�	�r�Xē�a����2d���9�"�rc�4
�$%F8�-BPĆYG��M?�QJo@���!���*~K�����AN%�)��Zo���ʵ�B`��H����ʗyZ˲ӻ�K����ʸ{{���\>�=;��2y�q[b��� �����Z��!찣����r߽H�����ϋ+�b��nk���*�H�:0g���GN��_��0k�������B�]���ǽ@���P�����ɠ��5��s�J�R�"V^*�2
�/%��g~L��_sg�S0���q�|��v\�AϹ�!����l���j���K�ңLjfN�:���3�ރ'�n��s�_ɽ-�"����~���g�W��<�������?w���
�sHXH>��XD��췛>q17-y���4�;[̹6n���ճqO��c��_�$�?��B7Sgh���`Jp��KU=�c�3��y.�I �ٽT6�4�%��hY"�-df�����=�2j\�=>X!$�'#1��|D-�f��p��� ��'%�� !s;w��8�������>bFË3������8���c��
�z{Ǿtg�:$�0Uvlhap�	s�/����Ⱦ��,�՘�U0lkFL�'ug����J8��OX�W�Qy���D�܋�gĀ�qⱀge#� k������t{5��{�R��^_�X%{M`/R%f����^�6�(�t� ��p�
�?�of����DQL������i�Jh�۪W��~��ZLS������X�cf�Y��&|&՗��(��B�ZrQS$���f���-X͊j�k.%��9{2��?u�|���ZR�����-.e��U�W��Wk�{�/Dh74ʿn���e<&���_�Ϡb�oa�bF�@�ЮB�[�������e�T�����nB_Q���&�o��Fx�]��&�y��Bi�`4�;�hF�?@�޲��x}�}��� @�pS~��v&�Xź���`8�N;Ǿ�]�s�����eW�@����Ϯ$d���2��������6��FU�Ȋ�GvSm�W���3f����/X��.�A�:��`�o6�ϋv+��-9�;�[`)^��s"���<��j�AmЙ	�D�l�ޤ4@5��9�*Qa5���6!���6Wh��	7x�+B&a��hZai*Ė���; ��A�j�]`)�@m�0����5�,�]!�����~
8�nT-�������,uK�gb2n.���|BA%�P���Z�OgE����8�lQ��+ǔKg/��!�����]�GJ�Ŝ� ��p�)��t���dS5��@�(���V�W�$�5o͔��p@�MW�gG�6��t���ʴ@ ��G2���f�3v��ݴ�tn1�u_*�����%%�7�p�/ZQ>Ƒǿ�qv����z��f�#\�]Q�`���P�}��l�%}����!��AIu�K�^�HOJu����'Em\6ɒ�60���sI��6�ʲT��?,�Dý1_"
����M�IPPDp�f<H[��!�IK-K"�����ɟ���-)�sրW(Cz�t%w�F����::?��)pNQl�Kj���]+|�;�\��)���o�>t�?��c��PV��������S*@"!��ʼ�8E�}�ɲVYc�����v��P�_�!@��3 ���H�+$��,���5`��ɝM<��O��!X�w��yp�'��M(W/W�U��3��L3�vl$��U��TS��,��N�
 ��Bڋ�����򧿸J�#��/�ݢ���a��դe����O�Y�qx��z:3�R�,r�J���m�\_vh��#kUi����[a������R�~���=_C��kB^M��Ji0	+���<$��@}�dm�9��k�Yt��Z������9 `�8�߃^��i�a~�F���&lb��K��F�	w�gZ\��Ʋ��^/kD�����Xl�n"��Z²D �ŵ(2k����ў Բ��%�������|�����P��D���<i�Nx�������� �����t��D%s�u�S���ˍb�Ӊ�c�?���Q ����cI`����;��w��t�S��*)uT����a��"e!� ��3��^}�!�j@7z{ņع��PT �@�q��'-p���f~���M�6�ˍ�VB�P1�V��ʄ��;�b)��8�O�耓d����4�s0e�,ʤ���9�R�7~Il�}���=�t��-����{��Vx��-a��N 5�ɗ�8���� K/\�\!
�u�F9����x��YX�|݆��`�x�@j*ŗ(zV�	��D�TPN�7��X���2�ѽ1d�RxUٸߴ@�����LQ,qH8�E�r����b����CQ�˚M/�Ń�����>���,ڎ@�XQ�*ݷx�u[Q����M��Y��l�k�/:I���->^!��֔+����/��)3E�-�t�y  LÀY>r��B���N>�Y���YS^S^WO����#a�����X�{`��T#��>�;M�6��w�����7�W��jCU_��-2��[��Q����K�#6��_-��vV�΁��Å7B�zf�i�G�icMH���ܺ'�O}�ř���p�8+���wKу�ψ��jTU��F���ܪ4�}�f�M�BtK����K D0��K4$����'�_��זe�F>�����/������s�t�ՏF���S��|��WO;]>�Ǌ�+�V�g�1��:+��x���U�z��g¡YP���bFq�\�	���1��� �A*�:*�U�:"�_(B���9|�s�}!j9���G�7*Y�|��Fn���ZrW�@�<i�B�9�Xw�ee������&Y���8�A���\�_��B�?�4���4/44%���L߳�	�ߌZ�� �U�^r+Y6.=γ��
Pq[jB�s��5KP\��1��3s�V�h�p�� �LO"�j<�۷���a���q��n,3k�^q�}7�S�IR��������&�:�V��c�j��a?Ɲ�s>Q(��ڎ��^$�!:��� Ybơ-����*���3�����D�$��(!z,���g�k�����}��$�� �s�Pq���%Vc�? x��U�d��E=�� �-Ρ�;K���w2����mP,�[戎����(J�ᦆy�Nʌv+I�q��K�) y�@)<��|��x3G5_�'t�W1�#��n���QoZd�M���%��1T1��W;��_�� �zC��ˀ�Yـy��(�����'��rZ�{촊�D3;1���n_
�y��꣙������l;�������EK6ې{2���u���R�������jǻ���ć����O�a�{W:�!�����6A�»�<��ʹN{_�I�\Zm�^��e�N�L���_ll&d�3�7c�?X��A[���k���+X�v�8���L��2)��Z��4.���in�B3�U݉�l�g,^�gx�&���!�$���鳛�Zm0P	A$�� q��y�C���]���b�k5�u�=�B��hy����m��-=P .~~�w���v�h������Ѫ����t[u��S�˵�1�f+�-EG`ʘIN��:P���S��V��Vk�zG��?�%�����;'���X7D7�|i�	��U�j]Ub?�ς �_����-���o51�O�^Eljf��:��G�;�0x��fTG_���$=ԫQ#�6����Dq���M3�w�Km_�S�������@ݶ��U��rG���� 'h���}�Kb�6�]�ߔ$=�;�hT�g8L�ݵ���x`��@�txp��L��#�h�o�d}�o�¿�.�����yrH��j�P�ָ��zŶ��S�F�4=���;�Ƈ�s.P ���*��QI�}��(6��B�T
t���!�/�l�;T��K�]�*n*ÓtZ��`��nہ��D�*��I�J��iƵ��1��cv#�M��Aك��&d����|
6shJ�xW�S��Zq,�B?L2��
�UhV6`�nQQ���p"\��ďj���������q�ү�ę���ja2}"����hq�k��=c����rkk��*jyRO���|w9���/#��Y�B	�qI�
�Km�����Sco&���6�8C������Mm�2�J�j~��kH����ӎ���d�eW�A6Z%�XB�!��(���c�v�n�<�J.@K&�����b��m���e��y5��~x���q�U;�t��b%r�?�7L.��^�Oj
e�eC.l�Y�,<D�2�boq�Z���Ե\!h��0�P��Z�A.M=U����-�
;M�E6ԓn5o�!B$�"����n�y�F��]rx��#�wS�R`n��������_�-�jCj�a4���4���R���&��i���\�3 ����1�>�BZ�J��ޞG��k+r���}�h@�)��l���MƓ�Y�Y��t~4��[d�.a�:��휗i��ݫk2�_����F���"���*�drOD)�YI]蜟���y�u�@Co �N�@�G~��a N=0�g��SW����@g���w6�g'��P�[����?<�z$b��d�+��oa`��A
Cί���.!�6X�
1�<̄�Hu�A�{�0��ef�3�TvY�޹`?�S�(��	5�N.��z�NŚ��p�c���[�a�g�[�#����&��l�B�ݱR�)��dS�Sv�p�����ٍS��M�i��T�r����7��Ҋ�'�xl�L=�R�/
���\3�
�о����P�R�W�՜�YZ:IDx���B�1h^���d+1�Dr`I�=�Ķ��U���9�h�.���`�Heؽ���h"��`9��Bz����K	"�����B�����d~==EˆqV2�>ϫ�w�r`H�9D�l�D�;l� ��g��t��r��|DL�MQ�f^>�V�?�=�3qF��JD��������iZ�z��hy~�����Fiخ�T^���u`Y:�Y�#y<TC,�͎��G�p�$�.�ۤΔi%�ByhH�++�FD_J�i��j��C�)<hx�T�n��+��.���_�3�^��IU��HQ�wb�Ȟ�T���jg崔/�O�����#Oy�jߥ�y�hRQᎎ.��[���?�lߛ�^ ��ʵ�Z>ɟƣ'��i�z5��5+��"�@"�S$�����&�� �Y3Ѕ�l�f�D�lH���|���Q����IC�
�,��4'�����kO�Y�S��e�g}A�xM	����7�1����.�mH!�^��1�5{~�C��?�5Q���7J��/��=�9��o9���.���I�����*d����m��͑�	�7���������cu�\�Y:,y�n��{��ί��kD����8�ً/og�Z���u���������m�N�̈́����Ie��\a�$���7E{�*�}K�K ߓd�K�n���`�vT��j5%��՚^�<P�f2�G�
�yr~���v\��mo��W����A�\"�oA�.�B�!�i�q]���'��9XJ�hP�Ur�yL��9ｭ��E��"t��0�;m�-tc��K�fߜ�PG�	`y�����؊�oA��:�)��D�I�?�"'S=�k�����G*��Ł3:ĝ��X�Q��K��R��s���>9K��_j��#͢Q�t��q���@K�0B�Px���ƛ�� $ �����F��z�	���x&��:<h�4�&L��U��l����Ea#a�w7l4H߂Ys��dpڀk9CD=��LqI9�Ūq61`�oG��a���[�����3��������ma��%t�n�D'C��b���)���h�(����v�t��oWl]���9gɛ��wf.-�_�;(���11hJ�YI�a�#��R�����_0	�۔3mI��O��`�h`���*���;:P�)!���zŁ�k3�����Gz�l��]Ztp���'�35�[�s�1����R&��n�|M	�L�y��1�Pd�㌑z���1�  ^��$5�M|a[���.�o`�\��O\u>q�oug�kE�OJ�e�3��7�����B9h���i��͍�n�eD ���C����en�7�&�:��Oϱ���Xk!(�5.���p<w��;�6t�Hv�(���>��7*�g�5'_h{��ӎX;n���C+�u=����	�5d(N
��_�zM�=�Egv�IZ�l7��rs�19�),�͂�`��("NuZ�j���6�w�D\oQ�j�H���,(3?|�)����D�z�}��L�p�D��7��Q�
�O�wƾ��/'Ц��)��>(����a��)*+��l���̃q+��S�?����&�t�Ky�O.�2�J����Z8g�{�\&�"�h -�( ˂H����ZNY�pF_e-��`��/j�x�+�u&m��[8nYtWB$Q���y7���E��Q( k���WYQ�)C��1@i��<�-�$����Y�%<�tx(���Զ_>��4��;w�]����aJ�Bd�k��Ϋ4.}���Hjǥ���V�1{n,�uw�ezPi��r��o^z ���UU�5�a�0Zݛ�*�`�B�r+��a�����>�]�_ �ssJ�D��]4�����>wDj���`�߹--~h��k�47ƫjH�$nU=
"����c:����ޘ_�*7|���@p�.&�}��	���udC��d�I����*5U���ݴ��c�RY��ҡ�*`�pW`
�%Sp�	F�^]>'ÔY��!H��c��@��&�w���a��}�E�=Q��Չa�Y��a��0߉�0U��ö�:Y�C���&�G6Z~<K��پ��x��&����snZ���#�u�M��EI��Ӈ��3���ԏ�J�e��yX��E�Jp��r�wyi��[�_�P�ZR�ږC�VDT[Dp/��%	���-dy8�R����B��/�1h�����<�L��]���(
�7��Y5�:�蘛��SEJ���f��?{e_�����e��
��G��HtF-�ΐ�g/?^���7�M�Bu��K�/���RrR���}���0�̵W�JwU�y���\���0��.��ʯ���헨�%���:������w`�������\�ݳ!����]��eDM���aA\���5���
��m`�XZm̶R�%\�����[�X�d�����h��9gC��:��j]��\��%`u�3��t�t��s�B��}�iM�tWU�c���.���^|�H���;V�%��9�&.%%Gw|X�=��`����H�8:��7�X��9m�pt��S�0l�����3�,��O��ׯ)ue�iPSy>ޢ��~��������|�?����u��;ي�P?�+�3�l�֘����)M�2��?cY�o�Yֽy$$=79�֊i�l($�:�����&����i�6��K@��{�z[�9��Ԇ+q�^�K��WZ��� ����:e����mf�=��D�˯�X�lhj�8[����d����A7�鑒׷Ra\�©	��o�K��Ȥu1l�?&Iz;nz��w����H�9��J�ݪ<�^��q���s.���J8"ׂ�gciV��;T�@��a9���'!���A��п�C��06	������m+��ȨJ@[kڒ�(	N�?T�#�^Ƭ�,tZ��k�k�~�e�
F�0?��Y'gv��b[���_�e}��6EK���W�uY��0ܿ��L���6��e�XC��$���gR��J�Ka/g�Z��f��˔��T�za�4�C@��-S'�ߋ��1���Р�	�$�@���.���p$&=� ��ǟ$�E�Oͤ�|��<�Ԛ{I����뤾T���5�q#���4�j7ꮂ`0��U�8s�@����mc��K﬩-�d��k��ZoNӛZ�I�!_�z8�B=[״焦O�ԑ��=)=(��ZPk�5r���st��Us�3�jo��f{#����z>�a��� ��n�>�sF���\`���ʢC�r��|N����X��!�uM3l�řU�C|l�)Zg�O�<.�I�9��ކj��Fc�#��&{�ƻ�i؅]6�2M"У�c�C+0~^@<��}����ƝV'�<P�NW�V�tԽU �J_�&��?z��x�M�|h�V�n�!���$ Փ@H�Nt|D�����ipz�x��q��P㙍�G�c��B���m�iwLX����Rg8�d�m����2fׯ+�eg���b
E|�{�\��o���)�-�4!3����s�>�ux~����F�"�~��4�W�W���Q�>��������F��a���:e~�S;�n)ێ���nl1V�A �u��D�� �S,jG|���ǃz�G��{����bbN�K{@�q���f=��m�L�%ө$5J��96��4��$�ױ�"ԗq��%�D_�U���|������oU�KZ��"�2�֧���v������[��d����O��ǐ/EP���N����_X����99upVN�1��Ӛ���� 3$�2����%���x�<%�9g�kv��GϿ��N�y|(��%�~^3�kw���pu���H��X��׃��o:��`c��Ml��'W%�M�Qy���U;�oI_Q��h��iJ%�~e��,w#�����X�����7�������M~S�K�td[KQ�9{�ƙpYx�.�H��n|�5��ET���7�T�d�������9��%%5�ס�(�*g���a�"K���4�LG\|�n���g*=�J�l��0��Tu�1���F�k`s.���1ձ�����Ո�Ǣ8e�_�ʵ���2���Q�'z��>�M���6�+M97����?;������e ���6�7�׈����z��ۓf��2ތ���������g�$	'�g�!���Цo"���@��6�_��7��|��O���	�` �W6w��@�8Hyz���F\�;���a��Oٮ�/]�pMۆ��ÿN�m���#`8
?"���������6>�
�^�ΤT��|W�I�+I9�4GI�|<�X[�@�^Ykь�Tk�
�X�zG��<����q�T�x�~a���[ǧJb���BmA[��I���8O��2� ���N�P������@R�;Z��K�Nf��O!���&��|��'(��\���!K��8B�7��9�s��F��=r�P'���W��>���A���RM����nm���5�l�&�~\����	������/ξ�W�MU��X�X��x��=�r� ���/h6p����;V�"���#���F=�������r=��N�������=~J�*���"�{q2Wﲦ-	1��r}dF��=�����[]�|��y##.��
�9�xӁh��p�`>-�H���<�vиU�1���!Q;���L���wch�*vX
[=5@("��~J�`�I�o�-�6�aW��F���u��E��C'�p����}ow?@TƉ|C7�E���b�~~ͫL��j�Ǜ�\r:H���E�T�`����������E�TD�O�����$�,�9h���3�:�W�]U����K��%8�<ό�c���|�����Ю�Q��併%?�����L���6�p�]r��k��H��y&0��Vr�$Я�`�}k�	+��a9SH3n�ZTÑ��o�A����l%Ӵ���K4�Y.:~x��̔`��{ ���}�S����F��S��n*xЈ��S#P���[�hG��ɵn��ɍ%���_λ���I�b��?��
�
r*E1�������BqZ�U�w12���%� �3{��^���Al������Z^��K�'m(3�R���h!�R�k��ü�	�JჃ\"�_���@1��n����.<��ti�I;}���7Ǚ��B�fYU&Ά�z��!��:�w+_K�=M�dz��M̭a�����B�]~eVgc�`�*���4���]-^���ϻ�J䜠�)G(}1%����@�yX��"�@1�QF*����C<����!�#k�{���8`�1*T2��""#y\�\bZBݪ��e����\VE<�t��{^���-\�trI�4D�\RՔ�I�̺�t<��O����7ު�{/Bw�9
b���o_fb�R������pg�.oZ[�����ў7�!��V�>�϶{,�+�����ڢ%�}ڗ�%�QZ�D���_�=�����רE���29��7���vF@[�Ր A�܊Oeplb^�s-g���4�{2�,�����~�����c��n6	R��d�S�W�م+�v4d�x �i?d��@�=�	��
�� e��A~ͨ՛PH�屁�nQ�4��L4���Qڍ{��g�g�$�'��6���h�۾=���u�׬x���3����CSK��z?��P��נ�����_�[#Be5
Ϋ����������|*ע?�$B1�������H�8vOс���6�����hq���q7��C���@^�͸�����d�<�a���ߎ�D��XǷ�6��x�T���UB3��~�=Ӡ�daPD���Л:�9�Yo��}�Rbb�U����&�5��Xl�ʸ��"�BM Pyl*���[jǠ��Gx���H���<��s�CK�5U�U�SOM\?���X+�r�� ������@k��l��f�/���2�Z�8>.C��������-��v;�Ջ�M�]N��G���SyWe����=��/���*��Eoy����R^��K=�nS��Ed�ѐ��:�#�G��΍��E��W^RP�Ir㇍�%�±�j�*d��H��*�Qag������T��v��}gx�l.�;����9ɢ�]���4%��pN�u�(t�����_���E��.����"���]��+�)J������$�G���y�ː��WX��5'�}Qo��p�)��?��ޔ	y�~j�p�z�ߺx�9�m��L,�(�Î�x3ae)P�H.��~!�K8�{dh�y���IE��d������P������=�*O�����Ը��6W��փ�0�ih�LR�eI�!k*���X�\��ߠ|��KDR$R�+#_8����_ar!��N �,M�fU��+X�\B�}Dq���j.�p"��6ح�ri[_M�S���*z�{����|���F�b��d��:����Ɋ"�L����
b��������DF�m�p�W��p�G��{@C/1!4n�mÜ��3��%�BB������@���:U&��X��
��!���c�����A�>W�w��^�a�G[��ݤ�F�;C!�������=��QE5>�o��|y>�ϵ;E-�zv�9���W�J��X{OZF�DVsZ���J~2��~Zvv���l�m�j_�;6���&�an��U��띋K�^�촞:"�u���z���aE����-����B��!}���D��R��X������Q�����I߻WO7<9�%�C��d\, ������n�j�t��������:��EL�֯�T�=��	h�)��&���R��I	ځ�c�.����Iκ���0�f���A�#8�TP�U�@w�Ԝ��i�Q��Sy�y�2-���o0���*WO��$��#jЎ(l����%|�M�^�*PK\p���k	u~ˡ�-��Q ^$v�)[���Xt�"�7� D��j�d�Z��z0��QF��oW�.ic7w7�9[��jď ^=QaY欞����5f����T��M��&��#A&%`w�5����18�Y8�fȭ�*8t�5����p[P��ɝ|����:�,tT����1{�ٴ����1S-��IR�Bi�
ʪ `��0��p�;$x�,Ӳڳ��J�s�oO����q=��Q�5����@]��Z`�ޙ ԯ�{� 6(GJX똿�n�⾎G�17P \�z�$^� c+?S��˟G>���f�%p�6:�V>!5L���Q;��g���(2���������g_h��ɬ��].�C����&!�7t"�d�z*�����J���F,Ք��Q+���y��4/�ΑI=<}aѓҳ���l�Z	�>ZI�R�&��^�^>�"ݬ3 �pɷ7if���y��]� e�~?z��?����P�:6E���>��(�ά��["�AY����F(��>> ��U;�K����QpGsl7���yHZ���}�D�|l�}˓�(���������_�`�zpJO�l4f_,[�����!T0�R��eތ����	i�B5w�y'�PL�Qj����m �ik#�}L�!��1�����H ��O}��n�~K>pи�٢y'���<�`x�L���E9`ܒ��FƢ�N�G<K^���E!$Go��W���+��(�P�u`��E�]��A{7%+0�H�Ӯ0�>����=Q§`4{���D��&�.�M@+H�G��{HU�U;�`��ְ�u��G���Xl�5c�R-l�P��p[�i銽���af��+���<��"t8ɛ|8�$���G6�yA��I�.��fO�s��S?'�jc�(m�b7�ZPeZi���9C�xy���n;�OO��V
��@�V��(WHT_��y�~c+�T�k����Δމg̵��gk��q� K�\S�N�-|��8W-;�/��U���� ����)�2��Rm�co��τ�Y�~�]��g�i4��!���"tsC��<kBQ���:�U�o��$�5@�Ү�+0d��m�iF@R��i1G�
���R;�����j�#]�	�
gKA{�zܦ�#�k��"���P��{����b�g�zU��C�R����\�<���� g�� ��g���u{y�忿U<
�?���7��9K,y槚��DG8̐G��?/�һz���Eƻ�HV+`�k�`\L����t�!�.�¢��훾��� ���\O�y��$KB�����4¿�:�j��P�[����u�����m���>�s}y-�y��3]��R��U�d�������δ��OmO.� u���^�Z
a%h��~�¸ٕ�?v�I�uaT�}ɗ�ONW�껰_�1x��X���Hto��K��F��U�{UPk���
�>�o�[C�`J<W�!qh�䁇�Շ|G#Mԝ��� ������s5��r�@��"_3>�����y��	h�;��]_���?/�8�*%=Me˚�t���$�Wj�Y��@ +|�tr"�7LBaT��|2(U-��G ��"�@��]~���),7D'�\�A9V�l����sq�改��`�QRK�af�������2R�-O�aW�>�В��hl8�}Xe?p�˯�G��,J:�>��%N�m�����=0�`�ߙ�9:7PəN��8��C;�(\�n�3�vA���c��=+r�Z�0$�x6���ǳ�dȕ���h�E���ԯ�z�_��'��%{�_����k&���,/��v�f@<���o�����2�o9Ƅ�?	d�;����k�BAkbj�`�����vl��|�Jt�<y~U�Q�]�Cm�;�{Ԝi�Pق;��c�\��K��~2�{���A�\oo0zP����'�P̶8g���dQ=�*��������	s�fe���v��NY'8���g(�"��ɵ'Q���> ):>�du
Vs���i�C�nt�P�ot���{��;�2�G��ȲZi��km�"��2����(�xJ���g��v�Z�JҀ��sL_@��'��ɻ���&�gt�O�\�Dj�Q�ii7�r���6���{A��)M�=�tu�� :��o��G�CW��W]��>`���ݸ�Z�F��|FRcj��\��+�A�DKZ����"�(��Q�ŋ\E��g�a�a`�i��=a��1��տ.q���ay��:�t�kj6��Dc�*�)&)���7$bM�8TJ�\�c�,���y(� �?��2|��^f�/���J��2�8��UIqm�8͊1%ً�z�+��28���M�X�8Pd����w0��Q�������/�Ⱦf�Ŵ�����7�v�0�-D�V5gnĊ�I.�����T�$�˱+�R��`]n�ǅ�ts���(�PP��&��H�d�]*.�� k�V���͈�sf�ύ�n��Qߓ��鈇%9>����"�;t�5�W�JC�͛��#�.��
E�uWQ͂����(uroE�ydߥ?�N�3K�ѫ��%4	�x%n�*�`(�t*xc���T-]��F�Yp/iN��'��W� t6�źK�-��d^w`�ܙ�sDJ|������F�5ʰB�	=�?�nZ��#!�ĪN�g��� 8f=D�haJ1+�w��t�ɘ�,t�'퍢�x9������P�t
]�I>���ۻ��r��D��cީ@�E�RB�ڐ�t�a�P��	`t8�¶��=ۋ�7�o�+4���E��j�"��\�Ѫl[#ٶ�F#<��0��F-w����b�R�YB���N�$����DA�6M�k1���3�<�RoӼ�kD<f>`Fv�|�h�!쮉�Z	7�߱b��HW�:\mmɫ��}����w1�I|B�f�^3�}ِ��qL�?&�Џ���	�8	�6�g0][n�Q�o\���}Yv��Z?KƠv�C�!�^�5@@F���=:�E��(��NB���a�O�Z����Z;L�'4Gl(b��Hӝ�EQNq����'���9��Vh|X�},������6zc����E��F��w�n�;�ꂸ�ܾ��������r-����	����7��*���mm쳳#x[8*pU.9�7'wox�v!�YeV^ڑ�6)D�`�#�=z#�0׎�n�@�`�N��y�!:#�������^�0����ڣm�Od�K��A��8��j�ƴ�_D|�*�h�qk�
���:��`hE�����k�VW�bR2J��q[
�~���G;��f�/��~˃�7���F���r�
��u������Xof&V���/ۓ�oS.C~�eJ����N� �����[e��9j�1bkDC����s$���X}A��"���
�TR�ʈU�
��/y�������l��,���5� �ԝ��10�C�<���k�*u�jV?��O�F�8�C��bh��
P_p���M=��յ�pZ,�Ú�fB�:��Ɉ�qV�eб�}8��~kI���u5$��+�/M�9�Ͽ�=�ް-���L�&���'����޷����,ZY����<��xH>�X�8SWr/��q�vc����e�J�D>�k����+X��Mk���z_$�xƋ��n���{�d�'B��4�*���5�<ٓ�-//�$lU4<(��&���8�^)wVgW�;OX/��C4z�Va��3���Xc���SKX7�o���(|�|˟������+��psR,��כ(!�1�:BgY����?�&�o��Y�cI'ZT��ț~�����X[�Q	�b�PV	�*�"�&�ܑ�wˠõjg0Κ��Z��d����3pl�9����~ۦw�V�Z���^�RqrнW5�W��1�Sz��F9�"�<�������5�Y�Y���Ky 2���Q꧶�$�N���l�H��:�o�)Ԝ;�rx���)�s
�W�}]�K�z������s=�x���B/w�ܺ<T�h�ƹ�}-��e�=wM�����)���&E�he�`�1�n �5a������eH!�Tȣ�-ܶ6�ĥ9a@���?�R�r���'�1D��q�.���mm5!'��`R�K`޻%9�,��j_I��~ �kwvr��4X�o�b�HV�b�����:���B���elZ	"��O�Z�]��Դ�����<��v?�ٮP-O�D�=)�+���q���|\h�� :2������j������?ָ�W�`��h
7e֖4�o~�Ƈ�"P,���u���Ȃ�]c"�N�EdU�&�~ل�GX)��� ��|Ņ��9Mr�I�s+xL��p.v$�"�s絏�`M���-X��Y��Ag��.��TVAYO.ߑzӇ%=r�?ѥ�d�	��<�7^����& |If�3�8?�n�[��YOZ��=�%�8�#��F3�N���Lo�M���q��v}ͫ�.l�Ɩ�8��6�M�.�~a�ΥF"ъ?���w}b�"�}�h8Y��n9ﹿ�d3J3�)2.q(��'�f;�g@��P��m0
����*t`�'�Y9;1����o$ᩦ������Ad~,��:� ���JqDf���l^�؁���
l_�7e�#��9�Ӱ�n]y7��+ȑO��=YUԼ�gZ�tDR�ӓk�x��S{����鮈�O�Xt������I�Ȭ�����6���yn��,�C���N�t���A�-�ܫ[��7����>����Y�6`i4����I�%9S�i/��:��m�����謖�Ҍ#49$�j�����lߖX��J;oq-��EJp��͘�xvd�O��uJ�s��}J��l�Z��J�l�_Is�֌��Ga "Y���/=���������ʃ���l�v��,��z+�v��O�q`�;Ja{�&x�Q��mJE1L����$+7`ۧo�Q?��ݏu[��p ɋ)���x�� ��� �0��J�t8�3«?ڠ����}i�WΕ�b��_��O1f{G�iL���z��D:�-~jm��n^�!�Y ��A�羙��1���˚Ț���
�pi�9s���C�
JSf9����G�/�}�T�Q}�V�SxcJ�1�o--��B���C��c��*����Ԃ�]4jF����
h���/���������+YC;��8P��6D�p�s�l�4$ߝ@	ʳ
�0ۼ��t����v1=�ի{�qY�� ~���w1B,!�)�x������������S��[oR�T���C_���� �t��?NZ��#%q����{��ԇa���9L��wT�g>����:Ug���]S��t��Q*8�����Z��j���� <T����$V3
)��)7h8݀U=RT:V=$�=j{��1pġ,�<Si(1ŀ+jTq-��9.둞ɐD'f�vI*�?V9��2���/ $�LV���Υ^���Ȉ-������ ?�g���.�:\���=�
5�fz�)�_qu�tu�{L�e���H�Q1����ꥢ���H�� 3�(�rfW�TcEh�T����R����Oj^egl�֋�� 	68�{��p�V'�H$��3���@_8���b�/
.)<u���EK�_����2E����]��4S����#��1��B���$u�Xswh�����Կ�-.�@�er�C{�QٽV_Pj�e�-�Hw9���a�"en���&�JfP?MJ}͹r�._JM�R ��*�ּݼ ���˟��N�?�R+��+ؤΤ=�R��H�����cde��	�Y�X��^��<���S($�����#/_�%���W޺�$��!��j�\ܬ,��8��}����z�ۘYN-�,�rLZ�R��gX�]�j)�՝W8P\"�(�*C�GN� _�
+�}i��) I|r�bW,|~Oė�/����G���g��.x�y1g]S[_�v\p	!`R�7n' ɒ<y���H��{�k�c��x�Y©dA�v�v��؜����)�q`��r��i���ds�jZ��p1.V_��AH�A�ɵ́[��7.R��&jQX�|��^�g������6Y�1׷�_Yzp`C4��g�P��U�_��u�K��m��9�m�f�Ѥf�ѐ5���b{�g�^�6����;G��*�|�H��r��Ŀ��fp�)����
�^�6����!���q,\�y7���F�N���:8V);�K�&b��A�
�:�2��.u&�sIj6v�Z��b0J~���_���_�^�F�3�JS�v�e�0��Mlm����/�8k�������t�7l�eU�Іɰ�G�E������P�����S�<�>(4y�*��(k�@�ԁן��k���kod\r(�/~�0��]�(H`�-�͌�:1s�ك��p�A�ěfM�������v�K��
Su2�8�*�~�!�q���)�(D�o���܂L�� E͉~;����k�WP�����jOƌI=0�}T ���f=�BWb��N�}�vx�^�PJ_��WG�ӎW2�#4P;�Nī���ێwp6���C��ׇV�X]��(v%!<��Hpk]<o�n����p`�e���mO�ұ����C���p#�ofOp!�i�&�p��XIy�A�Ym�0!WK�YS�\��=^wJ.dC1�����PY�h�W�2��!f���ϱ�'�JW.ډ�3�Yj�@�Z�@Z��ѐ~P��6?t5��ݶ�C5��Ĵ��mqz@s�'}Z@��e� �]GM�.1#�ՙ��i�Ў�Gr&�� �<�ؕ��~g��݁ ��BV��u�ld�p�Ѿ�[�{i@��q!������OM�����ɔh�H���ݔ�>�NH/�uD�(P�-!!`���p|VPH1�B�Fv��5���t.�IN��(�e
y^;�.�@A��p�lZ��_�P.�n�cأc��e[�M��깆O��u���YL����^�3��x'�����(�i?�J����֋&a�����X�(�-!Mz�s��F&�����_AR-p,[T��Y��`�>"��sZ7��s���(/EP�	���<�����t`+��J����鎘�W�A�nFOص�dVَ�j���<�+qU���E���` ��YJ?xz�����_q8M��I���.p���,R��ub<��)o\��Q��q���X��:�������0�G�q�c�(�8���r4�w�zĦ{n��1A%+a,<��T��"��n�G4��������S���`6��� i�7д�1��IW3&��ڑ��Nvy�W����1�����3]�V�MB��sAvʰ9����]9��bT��,֩��hO�U<�(B��Lgg�xԷsfPMUo(4�D~��9��ZWO�r]:ErD����0�"R��e�]��ʳ��O�-��7Co��i��-�X�'���}�sM�R��a��9�h�-	�j%�E�xo�۱l�����7	��<,#�B*��嗔S����?�'cjL���3�h[�0�@F��7/���q��S!��������* ��"kJ%��vF�2[��$�Rb �?Ӫ؂�I.Eq'[��8��ƫ8&fxD� =��X�C8[�5�"�0��\q��4��	�;��F�	��#�?Ȼ�.��q��+~��Մ�o�t�[�!' �M+���
O���*[҃�#m����F�=��s\)v�M��НY�V�;�f�ݨ�򻑉���z�d�RH	^<��u�<�ʾ�kK�CuEѯ�����e�\���j�@��
��Ө��(�~
�x��aF��L`I,�n�M�[s���AU>@s�d����h����}݊�E��)����E{3'	��jv{s��]�J����b��@�;�A�DViE5կae�		��+	&��)Ji�3�����ɺ"�(���Lf.��VS�m�LI��s0�/�Q�_��0]�d|Qi�p�=S�y�S��-I��G a��v8��fz����?B��N�If����p�?����K/�����+�PBr9Y����-�u�����r�O:�+ƪf�EuF�j�U�lĪ9�6	V5T�S���ӛ�69�ZW���[�~�)�g+��`�!�}�kYt]M��b9F�{�:f���zg����HO��.@�zgځ����Y�Q/�l7?g�̳w���9�c���Z�(m�N;�6��np�G�I������@�.�1��m�R¾�����ؒ�Kk9� S�T�ץg�u��\��g��&I��D��"�-ɟbܷ+�����j����d5��P�Գ�\�f ��V�PB�jn,ysR����Hl��P[
y�_�����U\o�lPa��p
*��~�=t����8=Pǰ6XCQ�[�w����iŭ1����2FmswG�q_��AN����΄Hƽ���Ӊ���-�sEu�P�~����Ij��wCp�����u*�e<�_�W�� J�i��e��m[A�p5	���~���L�PA�����w���G��g��k��S�Ex�|��9�<�C�{��\�&�����gA�O�G��=��E�]�u�J_Z�)�����%_��3c4����p���[f"r��E`;2ss�������)ɷ`c/P%3���_и��r_��Y�V���Ĥ<�ْ�B��c�e0w�4
���˩��oKm�!�}��N��2=����Vզ��f��x��j{Eo�ڽ]�qlml�ʷ��?@?�܌��u��D�(������<��ɕ�6.磏���k|d���!:ZӋ�Z?�\�{/~ۻ���d쑛\��ty�a��P:���X��yG$�uvĄQi�厛�:��M;Io�%����(ʑ�K��U�~f��ZR���"�>�U�r��S �c��|��;�W�þ���ʷ���WL�(̥l�KH[t���uYHF��o+vw�!V!G�D_Z�M��c�`Z�̽��p�����!o�����$s~�<�����!N�6z��PG�KR�a��s$/3N�g;o�{"���HR�es��֑�����X�����P@�����]�>}"bW���z��i�f!�{G�}�X*�8���b�h�xL�X����{T?��g�u2�5ќ��\�c;�+Jj��atz����t@Ю���o\�+Õ��J�?�yh�%�lT�FPx�VmX�����3z�<�]�>o@�=���7:�9�{���K���`#��n���i�FI4�2,aN��r�R��-��%�dP$�<J�P�YC��ˑ}�.%�mE�(���G�Vz��L8�Pi�y +'iO>�T��h]?_�М��)@}r��A[�ԹV����@��TLQ� ��2��:g�4������[�w�ue�{^y7�t��[ u]��{�x��{޻�e&fF�D��Rm�ڔ���@�@�ĺ��3��~D �;�lE�1��ˇ��ɹ�SryO���5�\��ʒQ��cy���ԣ�˘i��Św��¯(�T���z�Yu�n����074���X���C���.���pm=��Kz������&6����xkX�@���Җ�83L=��=ME*͘%��m��J��H�sB�<����3�u�62b��Üx�E޽�$fgD�<0�'��d���0��&�3����x#ʍ(�+���䍁NN'պ�����Q/�D�^�2��Q�o��E��t�����2k���2��S�cښhR���3V[Պ�d��'���C�
ܞWoa���6�����p*�ǿrY�#L܅OS��}Q�i@N9��Ԕ�]$-E;�Fk��w�`��wn���z@j�������l�1`m7�[�������y��c���N���'2юU�f�d��ܬ���7�~f���x��MA�yV�d�aY�0�_���mnyMi'+����N-��vj��{��mt v5V���L�k��݋��I�̆�+���9���q4�(qW��~��s*���>�9q��ذ�Kz�73:VPtY���R�_i� [�
�/Ț �䍚pz�9�(� ���_�">��W�zb���������L�SC���sM烢�a�&��GB��ǘ:��\�X3�
��O(Pnt���7�׬,��Y�!?���~��$P7��7�.E�k�$:�Ȝ?LͪD_�PZ����}�&���s8��,c����1]�&LylW"��� I�ڥ�?|1qX2��� �H;v�_gWh4��Hxb����Jˋ�m
BҦl��Y��aben�`d���}{�)�jؓ�{=]�3�bϬ��)!�B��}hZ@P���u�~�C�2��7�L����~�7�W<��[�!�>p[ A�N�7V�Gw6y�����u\�	�b�Ր�Z���H�܏�+�xT0xK��٬����/�oy���22��6��=��qI���>���� �2��,��N�����6�Hn����Dc�mhY�\߂+�2���AM��z�����S�4�g��[��
}+Ի���Iv�$�)8�@ ����6�/�d�rB����n�6{|��U6w����W��o����!݋��Y�Ӝd���J�v�+�,�8�ͤN�z�m����I�Q�&V���=SX������/O���c��;��u�C�5���I?�z��!�h�P ���(�ѳ��lk�l	gߞ�jETF:������(y&K֔����%i�۬��UD:�٧v^J��R�WG��ُ$�ƀ+Q���q��4ǰ*�� p5E˰�@z�6�&ɱ4��M��$�9v4�o)�1�-#�/t`�WX�Br�,�w�b�����Y�or#��	���<�Eu0[��Emg#SP�_},���Q^���H!5g���;+�́8׌�~���/.��d��m�q�:��3����Ji>!W�̉a��m�&U�@cj+��M��~2>
3��'@>F���X�?�A%(r�y���S�e�.4�		:W]�)'0V�6�⤭���$=Ro�u�v���u½��2�Gc��Ql��#��iO��|?���j�Y��_!)&�(*2:2<݅p��]����>�๰`ב#���N��K���7'�{�WA^X<�R�˦�r����d�*�����@[��䅪�~�@
�
�ɾ{|�x6�3w�E�����;dSX2+�2���
�ZRN��eI,����o���0i�;ڥ�$;Z��{�oe�JK�[�`������#I��Gj�ٵ���op�A�
qZbեH��<i�ޚnK�Ye��ذ̓â�������?Z��;�w�+,��j(ؔL3���&'���e`�����97�d�V=�����8<�Nl��S��k/P�e���K�@Jn�S�Iз���&�Ζ�@]:�P,��_�c��)|ͩ�تY�yvrk�4���̘��Nk����tF
E ������S�Y��� �}��R�j�_���P��$�x��7	��.G��!�,�ˌ��~����ò{�N�%vw"n���m5��α~e	M�Jz����:��V*p��֤{[��E��e۶/�lV�� i2�?�7/�謍��umM&��]bǕ�_q�[[F�������~�D�����"�>lI���|Ʈa�/���zҒ�3�퇇l�r�WV��e�ϭ��w��q`�������̛�.B��[�Gm,�&�)�6�g@RH�ち�#yF!�3���,���0�{p6{�D���O�-��o�zEO���
�gKq��Ae��`���:v��I�:��0���7�d}cͰ�:�(f�I�V����Xz�M�L�hB3�W�f�zM_Nt���q"��x�]��N�ΦAV�~� ���pF���ʩ'�uY����.݂������s~��b@W|�X9/Mc��1�g�w85!�s�S�i,%%a�X��p#�*a������M�{>QN<�������,&�^���#>gv	3R`|E��	T�{�A�@�/Ud���p�%`M_�O��Y��A�We�KTU��A�bFz�WU)��Z�k� х
�������3|�8k�Ǌ�"��<���"��Z�pi�M��#}��7m��E��>ܟ.\h
�g���� 4���d��</�C�>�����)&�b��I%��Pkؐ�X_��8�N[�)����M�W	u�x�z�@�\�I�#nE���-%8�U��;�c�������P=Vր�]�sp�`�"5ɫ+�\�$/i0 8a�1v���ȡ� X��d���w��M���c~����Ji*��?�
�e\����	�$C`��b�;>������&<`�j�w@��b�*0��w[�怳2,�ް�^(��+8"W�n�K�(�ڟvڽ��{����,e�y� �1�����t� 6���,+���"�����@gɫ��z,U�Q����+�R}����%����:���^�/�Z�p��<��-?�m�Π�]��Iu~�yX��[���^֦��?�g�秩�����ӗ�8�/�4>�3zϡ˙7��V ����kE�l&��Y�})��<�*�Tw�Eq&�&h����w_Ѕ+ZnR�������=�����AD� ���A'fX�y����H�g��a���KH>a�٢'�̿9p~�[[����0���?�I������8��PոS�!!A�Y�!�7�����ȱ;�6<7���>h�X]7.+�:���Z�lө�RB����M�����a�m����{蟞2�d��+���~�,D���c��:�����^lF�3�}�ȗ�����~*�\���=E%��9s,�5~tˏ����р
6�U�ڥ?�}�v9C=��1��Y��Ӳ'�s���U\Nךt���hjK������1���m�!h��5�C�:*�K�<%I������I�@�� x�	��L��Ce���NW��]I�R�*7u�<��u���?Z�[�f0ǧ,)Ð���V6�RT���I��y�sK��c�%�n*��-����������Do���"�k���E�4��x��o�y�R|��9F���x��;y��G$cc�C H/1IHX�yҹ�Q�(�6$Du>ϱ�
��;c6n#�P��N��b�Т%N�'5�|�ei�Re$S� ��DqQZɮ�t�Q�w,Jy����6�Kp
�6�:��x���t4\��ܴBM�m��
Ǯ�{�*WxO�E���"E�.JI��"�RDyS��Hً��CT��d^cT����)���lRǣE��nA6Ӈ��ڎϣ���#�F��\	�X�I�@��ʆ�����QM�3=�;�#�醺T)A��)���>Tz�yэ'Y�B�x�4�]��B,K<w�sJW��Z,9T�@��̻�������?����>n�D�r��9�bX�9|";q���|P\Г�MS屬~z{FvR��%|D�$��� NH�"t����(�
�<�ʯng=T^s�i6�@m·[u	�(ｵ�3fW�
��W���9͏j��^t�"���UJ��y�-�DY7��"��>Ҋ&�_��4�����I�C���ӎ�5H����6@�&_u����~�	MPB���4Ύ׷�7��v�M�g����~�����c�c�Y{ҏ{�<�Bb�L�����ס�(m�ol�o�Y����Ade1�PhV9�k��D��邙d�c�9!�y��i?��a��)��� �r�mU���qL��<�g*Hp�x�Ћ�`��C�f����3�X�u�:����lB�8f�^�?߄��%�Yۃ��o+�w���l�o_}�]T�f
��Ƽ�W���0�ΡKDJ�q^5�F~�ԋ��=�a�(�'� [Ȝ����xtATG�7�ף�H�9>�a���TnVO�d����4�v�_y�����K�Q Lw��d�+OM�+N�U_����bd�$-�K���dT,.M-*���bJ�w���|.݁��?��~�m��k���i�A9kL����^IV8��m��:��n�̍ �/{BH>�k�@M)N��տ}ج!"	}e���]7{�.		���{�-�/v'DVP�m�jlX��:��xE 1׽E*/�g�7�����~��1�x[�b �3o���$���F���7؏��CG=�)���U��> ��1~�R�"6��װ\��n�S!&,����t�%��S���m`h���:�.<����>�.��y��z����5 ����`�9�1��>!�I`�,��{�Y_����d�,�w��I"�:��4����p�e"ZB)u��;� �@���2�*|E_41~V��`S��B�!8��y�ߨ�#-��Ɩ�1�T������&����<{����qKm��J)o�_z*4�qIa~hK�o|.�\����h#2P�̕u�a�[蔳�z�>���s5��) �G���dU��<�WW��`}�I[m��q��M�u�9��!�$�^B�`�����3$Oj���I}9�\Y�ڱ 3��@N �ɖ���I�Q�CqS`o�����6t�f�N@Sy��WW_�B�}��3`���f6^T� ���X.ٽ�z�Rٵ�]`�%O��dg@�2�9�K���F������q��������	���f�c���3W�k	֠�~���}ëԤb{*�c������Y�a�+5���1���Qtr@i��qj��-����JU����Ph;�&V2���,{�g
�iF�(O��Ǳ+�k�>�m-�����u�F�=�y���i���AZ�"�@0��!'[�ϣJ�XEb��J��]�4�q�L
	��C�V�=@��RK��Ί��wB:O��',�-�#>�j ����8�f��� �OA��k���6��؜��8u����5�(8�^G^���f�_�p��>|V٘����$\�2Ō�+��|
$n��e�wʼW��+;�[?�����owfD�(P�z�jW��y.����@��$kQN7���ڜ~u<d�
"��E 5�[��k�N��t�ƶc �9��� ,IJ��8|�>�^����:��l2�hך`>Ð;3d�����������߼��[cha�N8��]���NA0�Z�[��ihOl���d�s���=8�`�`q��Y)8`��q�W��숌��0����՚v����ֳ3��ʛU�ג�R?oqr��i\m3���0�Ĥe�c�zo.�x/H:�*��l�	D7lS��81��h�m� vo.��� f7ۻ��#Dk�
pmZ�NNH��@)o��}xyk>�T��zۖ����$I�	0�	����vw�ItYx}@z��e
����i�S��#F8�Z�da�ǒ�H���1���j=U����U�"DN�3L��
�s�6�3	����@�����SO��"\Kƣ����U�Џ���/[�M;̂ܖ�y]Rg�wX�&�E�ΛT�H�XM,-H>7�N~�1?=-$q���ʚ���|�_i;�x!�c����+r�����Jz�\��rc��n�Ι%�N�1�ϟN�%p���uG���QVvn�r%T��`��f?� �9��'V[k��A�{����{�AEoc��o��x0sc,5�Z��i%��������{������i�4�k�C����PK�4��"�=U�0�����X__ۛZ�a�����b_�-�q��9� �[�:�4�:ZzȎ�Kɓ���Cl���Z��p(�}o统*��������Rɩ�'7:/���J�,�w��C�@g�{ ,Z�hrYT
r�ę�E���+��,����h�łYX锝^�����j�)�/��TY�UfFE�?��Xr�2�rf�J@~��W�.����<���ubO��Vj�ӍT[�Y`x�����*PxE�����sAُ�ʟ%)�S?��zb-�D���xQbp��Pf�A�(�1����L��|��S����e�y�Tь�
��z�w�߰'^�����V��`~���g�C�n XX!�����G4Ҷ�];�Op� X�?w~��6��,µ��Ũ�~����?S�CZ�l�,n����	�b��ʌTVk,sv��ҳ�;��������?�'�Z6���NZ�$;*����"f��~�擽�j ��2Zh.��
W։����߻ 7s:���ܫ��JPR�-�c�PDHӸ���� ���x2���mcu���m�����O	���ĔZ����9�2pB5��>ov3�թ���y/of"Z�/�}r���">,��~��#���^�U��c�?]ԧh670�66���ˣ�����)
��/�)�?�P�{�Lk��TR��,��u5�(�?y�O�1��6�9��!�uB)Z��H��8sL~��)��H3�"\��qc~׍���=W��1���{���|)� ���5�F	x�7W��(��V@�m�s"UrbI�jN�IÛ]�󡚢�(��1�r?	�����v�n�Ï�LLm�c�r�p���8�2H���h�NKvF��2���q�π�I��X�E4�C�R���pe�-3�f��0S5&�_�M}м�&S��nw��m4ܵ�@ݦ>��>���ژ��E�<��8h�ߴ�yRN�*~�p�}(� )A>(�p���@j>t�涸�9� �LWiip���/We����B�v�t�IgF���3���K+,g[�Ρ�����c-��E��f��J���
'n��N�=�Ț��r�Yʰ�%��x 8������B��\��|�K'�� ��>^K��t���X�i�I�|}z���Z����f�j�17e�c%����n�@��#Z�R�W�nDf'X���N��i�R���)o��7~�؊n�n����OU�4�+Y�I4E^��z�g�Sˣs�rʳl����L ����V�����.c�ج:����V�>�-F)�A%tG��1!��������P3��<�Y�!�%S=��#<��;�j�ơ�i�?]�<�61ЊJ�A4%;��3� ��e�4�����뢞#RO}�߯1m�� �b�M�㘄x�Lԃ�
���һ�_�Ѵ���D㨩d�[|s�V�_-�YS r}fo��o�k#�3���pj������rV�2�n&�cؓfpÂIK%�;/�_�F��eŷ]o8�v���Ã��s�=^�X�X�p�?�ؿU�_�1@�*��O���'�m>m�z����Y��o�p�xDE��SS����n�O�k҇�OP�Ϥ/�KW\7tx�ꆥ�Uv�p�h���Lv��~�+w�2��CD��i����R��_�q8Li4�@���D��LY+�~�䞥���N�;N������;�Ǿg��ʠ~�6�K,���R�5g��5�:c<ș|f>vO�rG<�4�0	0ͳ�ղ���j����`�OZ�Qb&uK^HNEߞ�dQí�$�@0Q%���2+����}�kA���Osh�׌��S��U�-��(�� ����g�D�,UF��0��x��q[E�Y�����`WfK��Z�!����i��P�()3�~�&F�/����	дX�ɠB;�wrfޱ)U���W�f>I����j�jƟ��n���3����Աm�a0�c}1��bH�~�A��=/���>�R�,3V�6-���L~
���^ب� �&�G/W.c�G���R���)�����'S�
(��H�]� *�|}FWtA8����k�܁\���=u[R�X��Mq�[КE�$�`����3�uE�#J�ޥm�~���\o�%��M7���S���V�A��*��H7��k���`A,���ݫ����ptV��?	�S+%%yo���v4�W����=����gQĮ dg��i����t�U%����R$�����.$��J�6���IeG���Қ�SZ6LK�-m�]R?:�9����_'4Gq_��8����c�E9�-"RxQ�IqDO�5ìR�V������1� ��\G��ꬪ�g-�qJ�U��p�"l��H$�F���#�������=�� 2�%��GpE��n:��O@5b�=�%�i"k�XmNNB�;"׌:�m5�b��v��ZG�i�vݟ})'���x�n�$�;`��غ;ɢ^ݻJL��os�!��ڙP�c��<G���l4;�đ�a��OAN���"i	�4s�M����]���>����S	)��SFtEE,�m6�Һ���(p~<���^aa�L�c+-�˛���r�9�ʶ��&��g�����a���R�o�7�L n�/��%tY�Q�ř�@Ώ���I��c"���C9��>�d��FH�_�� �^�_���pƃڼ�`l�6��[ro�sPT!�;<��4�m�Z{���f%V��^��������rA Z6��T�yN�L(z�V�+-��=���}��������qZZ��CKT��x���Jt��.}��^r�d����C+�� C:���p?���4�=3=�ц>Dg}�?�=Ars`� �p6[*MQ+�¤��,��t�.m"Q�L�rG%��ܮ�\Y� ��g�/��0�@MRYU)�
[e��OV�p״���BH䨖%pYPa�%E���N{����_|�҈b~��x`�Qb�OA�0���r�܎	�w
�?��\ܻ@{�>!|�D�͗Wa��A���4~ɒ�y�jI\b�������F�k��"�C,�lB����P�N��o���g��&�D�HӄQ�p��ګ>��o^owp]Ӈ;9'z\J���\���D�闉�@����J�3�Z���9C8>����u�H�|���.dDf��&�KP%�2̮�2��-y�IH�R�|�տXU�_��ln�i�$V�z5b��]�*w�a%Y�\��V��2�EEõ	W�.((�Z�p+����4��F{������W"��bD�-��$����%�ݓA����S�9P�u�" c����}�Ĥl�X�3�s=�: ��l@����be�d��\�Q�Y�5�Hi���C�>�����		�G��u:�4?�M����/�P��������v�0�}� �n�̆�4���]ӝ����Tq���}�j�-[�$��]�b�qwЛ��T#Ft)�h.VT�nҡ����9dV��ޚ��Ӽ w�54%� "6��_@g���x��mu�T�zȬ8V���N�l���)����ǚ8��(���k��,�T&N���h�=�<b����>��4�����EP�S�pW��̑�&�wm���%���ţB�� "���3�W��AN]L���Q-��򈲣�-����Vv@�Ғ���(��������p"�jX��+�I�Ia��C��6�y�9��O 3�z+Z���Jxt����FTf Tm�W�`�6� �lӰ8Ϲ������bv�s=�r3��V�7+�я�� IPM�e��H���]������� X�F�m��5�<�{g��;�1O��E%���|�JQvx�*���Ġ�.L���0�꯰�_yܷ�?Qj�Di�xz]�UM4îiܱ�s
>�O2�Axsdy��Z+^ ��eyMpy�{ڛL���gAv� 8xHyb΅�����K�<U�|�j7�,��"����*�#e��3�fZC˘������g6�'�_��>��_����1�J�����i����0xk�U��	���d[�����7�8|�2���So2��\����l��3`��<Pa8}�T��V�Z.�Q�~+hd9�LT������P�!٦+��_L}P'�j��ѸTh�j�ɶ����(;��N"M⑈����<B~��M<�{��KX�:Ev�;*Ѫ7P�pGp�/	���� 3.1���,89����:� ���)�!ө_����qE�6mr�Q�@L�^��W�X����:�FGįS$�n$�y�*e-g;�4x����Z3U�%nn����l��<���0q�@�●�sK�r_�_�.)��y�A%���\�L|��o\c��8��ɱ9��(�a�DB'ob�ǻB~����ҏc]^�zb��D���R=���ق��2j�{?S��C�B�̥v�e��k66F��	yp*�O�j�L>��ZO�18�r�NzKYއ�T ���I�|~�.3�a�������L<�����Z����V�
O�[�������U��lS�I¶ɀ���N��E��=��հ����h�&�n�@!�$J<��Ҝ��B`O�_�K��P���Z�B_G������1ڿL�X�8���q�rR�^)�ԭ����"��5�9�L����}K�Z��H��1��i�u�(J@��̶�Xt��+�[�Z�����xa��3��}��WypVڤ��F����-eT����C��RGi��4"��5Sۄ��D)n�IC��s,d�b��Y�z���֍D ���Sk��A�'Lb����[�{X���w@?��Հ~ޛ9�oŋ�E���*X���R��}�-���oiz}P�9#��F:�$2�_��=z/�tm��T�-�5����h��
���c��b9֞�)܌���F�=�6:��`C�EZ�&���7Al�!©h��-K�������# �vk�FC��z@��& ���6��"�J�p&*/Ϩg��KhE�W#؋���=m�)���-�ݑ7���n��F<z�D���T�b ��ƝL���;�~�Sl�_.�D9��l��@@�����r�g�.|�Q�y��^XB�1A��D��a��C�H��N�mׄ��NKA��0���)��8���-�Yk�z�)ڊ�ɥOZ2������!�an#(u`bğ��~ݡ�.�ڔ����;��{h�����#7����/��{d��kM��E@`LnCk��kt�3N��o[d�b�E��>�d����$�+����c����qM[�m֓���:j��0%�iE���a�Nֿ�v|�m�Ҹ1��|EPa����*�� ��~�Ư���\#��WO(���@����R8�#
���[�����[�I��x�i	�W,���_Zk�����w6H��$���.�El�G�m��EJ����̔��iy�����V�s���G��x��U�b�t��]�q|Ĥ���m1�P��F�S#U/LE�- ���e&a���)���Ȃ�~�(Lc����"��vؒ��N������r�#(T�^=�ѥ%���j�S.�Վ���G�Re�2��i+v6lc�B/�v.6���l�PB[{���- %�n5��������K`�&}qs]U;��̰�8b�
��р�TX�D��S�α�e��a����A�3[��몶�����p-�$���J�;9�xWuy�L*Y����LĀĲ��W�$g�h^�����-�' BA.��Ь�kyQk�Q�R������ह��~J�9����
��D,��ǅ }� p�"��]"+fW���:�Qlf���1�Î;������o��#�^Fni> ��M���t��dy��@��ŋ
'ߋ�L��H(=�T0�]�v���� �5*٦9����{_�3AS�kXҸ2� ��(u�Tw,��Q"��^�K��{>w15�M��#�a���Q:�� ܀��8�;xI����0�_��K��W�����蠡dc��i�>`�M��U��N�7�{�_kj�g�:.��͘�_�90[:+Z-�A	p!`X�Ƈڱ�9��[�(�=��I2����P�~??����mH{� u~x��q��9��+�]�<96�?�^�'9i���48v�J��_oe��pT��A_���n�e���T��af�Q�����">�SdCU���)*�Go��Ô�y ��:��=�?8�׾P���#��k�S-��|y]0��%n���� q0�\���썆��?��K��K�.�& ^9n~`��F�Fv�n��׉�R��!�$���#�Âe�[�t��%R��2/|�Mq�z+�GΖ�!��|S�N�T��>�YK7Ņ#p֑"5�AV��1�u��|�g52�;�q7��W��N��|��m�՜A<I�)������m�-�U
b���(W;�+���|sʜ5j#�$b����q%�ַRH��P�<ۢ�kf�#�?%��=3�3!�d���<2u&�}����]�:ˉ��T�1�����A��2��-I���دM�_������]mT��\f��T�]n!�]��������2��C��xX�y�j���$I�R,��2n+���|�iA��	���2�]��*�2����!?�U\:�r/��A:L3��8���u��H��u��>evjC{��;����;�H��Ÿ��nP���U�	���F�v�lm�`�J��x%�F�3k�?�R�=�}}v���̺y�����C��r���ߎR�P�Í�	���i�/d���a�@j���o4(�o����@a�Y�bCkmqI�A��tS�U�@��2�a�A��L$X��5���|^��l����}M��Hh�$k b�Gf�	��d%륆4� �C�?�7T�*@�]���Z��mSxŴ{M����?׹Aܸ].{�roY�(���3�����H�KÖ���[}�/��E��lW4й:i�B�2�E�hLO��Ez��g�\eD���Rѭ��#)�\�M�"�2{����k��nm3�<��b��'�f�X�Ie������v�xs����kD|ٖ�W9�E��8�gX��tw��'�~"�RŦ�6
����>��L�I�u[+�V�ٛXB�Ve@�y�7CMf?�%a0Ff��O?�ޮ�hO=3CF�/0��p����inq�3�}v"?XU�t������_�k�sEm���m4�RN:"������.	��&m�@�r�X�(������f,�?�عeL齀��.%S�qX�b�q�Qp�Y�+S�dk��Hԉ�+�-D�+�5�wϿW�d�\@�.X9�A��<;�U}�"4���0��c�Z�9X�t��*��8�3����� �Ƹ2v�������E�e>Q���U�K�F�J�UA�ߢ�5�O���_���0��+�Y�H�Ú����a�D�޾N��ks���X����F�@w��i�P�Q-�҃D���LƿUÇ�sLF���ն��?=��%�¶�:����@�qR��B��ҿ�9�ΉN��kE�RX*�pr���U����k��꧿0��?���[����C��0* ��i��y<���t������ �(A'�nS�i��\�f:v�R�_�an��ϔw�hU����U%�|�?=D�`��q��E!+M{�����.�o�G���A�����h��;5j֒#�8����rϸ��W�J5a�X�]���H��;[?.���m6�>���2�	��L��%��_א.������}H[b�s�6@�fjS\�Q�^�Au�k'�ߕ'ܐq���|��k�����K"���B�|^Pk�MaE�+d�:*$��$�@KjS����>a@�ҍU��8TS�����ټW�!Q�V�,V��ny�v���:�3l�\���K]ncA���7eF�XH�:v�,�M� b�H�Lψ���]#,!��_�������Us1ZQ�s$�Ip�����<g��*�)�g�3}q^���@[�tR�Á*���R�`�n���rd�P%!�x��0,��o�'π���?�ͼxH�g��1�<��0*���pb�]�|ތ*[@R����F����m��=�[�젵�f���{ˤ(3��+2���u<���_(r(��/Z��=c#:����@���'�2��Rz���1ԇ�CZ��y��ӻ�M֠��̖����r�Q��O9;�k��}ds{}hєQ�?MxS��˓zK1�tBE~��>CA�8�d�ٟ�"A���r� �=Z�N��W�����c�L��N��;7�:Qs#@����_9�i�h�yz6 Cf������>|\5Y.��8W��r~T�~�M��1�j���P��)<]~u�,޷�ꭔ1ީ��F?���F�����?�H/aY�H]rop��l)��*C�T��y�N�L����O�=6ղ5!��DjƺУ>l�P0�.���L}���*RB���w�L�D
��}h�Q�&�H��H��Uc�T��4����l��,h	λ�T�ƻ[�Ѵ�!�ٯ�_{�1W���Z'���FR #m���y��C��
AU
�C�o���19���tw��I!�Y�o/����y�䌜�����e^�z�o	h��á�	� ρgK�՛b\{X��?
��\����[��" �"7sB*�-ܘ7n񧪑.Wd>��e���ѐRi��igD&\`w����(�0���/��K��c`D�91/B������fK��������>S����]�J�lIa��>y'2��k�L���r�+�	�yFb�}y�+�����_�`�OJ�~�!��D�a}*}��W�WIVOp��`n*Wá�@aD���=ۍX���tGtl���8�+�wQ�����G�+\�W����Pd�*^��Z��8�	��n���������.4V?�?O��_�vS� �;��������g�1��@#��*�V��TF��h�=��>�(�3���iW�B�N���ޝBg:�=&��I9�~���wD�s�H�˭+K��v���8��gǀT�! .~�'�R�YZ��W�U5��A%��A������iuƦ�q�!7R~?C5�rH����n,{�_�I��kT`� �-�z*���t4���u�m�����I&���]��-b^L4¡em٦����"3 ���=\߉����9��zm��7E~|v9�`Hw�>�G��j
�Vn���(�	1+�G/�'�!�����,԰c����
�I��M����i���h�E�ސ�&v`ɼF�>3�_��6U}b�l��Arr��󧫢����%
���fS[&4���-�p=��d>���;Bve�&1�6!Z[;�v�,C�3�9cpt��Z�� �kC�V6cC��3kl$〨�筈����Bh���� ~��R���l
s�$�*��~�a�]I~ 5g�*�mSe����b0̋F�dP�u���pK��Y µ6�>�7f�O��%�lH�g�%3s7��_�RR"�����/mƌ��l�4N��έJ e1>���r),=Cǈw#e��Ql	�CϢ\<�۳>-�S$�댏�n�͙t��Iu����.�F��ٰæ�o��'��
����TJ�W{�:� >��`#�)P�$�C�����i�e���'��ЗA��H�9V]m�qp���뙒�g����L�#8��������Yl�|ɱ"����~�3��%�*t3�B�^�2פ��au�g�\��q���g=S���U��!�f���﬙D�ֶ���l�&?���#�����,c����;��)�n�}�n3�.,�A"&��+
1C����b����
���>�$IJg�忲�*jB�u�BF�I��OɆK�@�E���.mo���6��>�*����x�Jb���
��Aޮ�$�D�\��l����[%��f댕&)���8��;�&�8�h�:"B���D�`��甞����{��E8S����>�|�����5��]]DL�L�Q[ \�K��	����4�)疆�C��1�nr����d6p<R�'Ph��qZX�i̿�{cn`v�S�G���+�IF��:(��%�X��K��sٕ��߽��]4,�5�.j�1f�l��?�u� 
!����� Z>�(��
o ����<&�B�L���2R
�]�����.�k������$z�C*xE�FN�^�q�Вԡ�M#�*x���1��ܳW�~DK{��w��#��vG,����l�>���n��k�����U�<p	�TN��f���!� 0�cP�Tu�~�Pog"V2+&�n�<���6a����߅t	�Zˉ���-c�Di���,�q��(A#�Dkc�`��D��~�-0����/*(9�ԏ�Q�,���M<���q�ڂpu��~���ܔ��s2����w`���`4IBC�g4n{i\���G*-
���!a�"�1�*V�T>>x��>ݟT)t�}=Zl�A�=�Q
T�oK���ـmV�7����N4��!��B¹�-�t[vo {���%j������=ޝ�5�b����$�)���~-��#���c�Au)jU��� ��g���s3y��ꚱ6�*d��:��8��J:���2�G/�I3u���fF�����$�|ظ��ERn����zR��)L����R�&��d�c՞S^vPQA
�i3�̛�e~�eº��T	�4a�R:�I�t΃���)�e!-����q��J�1�q|�_`��J2��E�u5�o/��.�~ݫH]H��!��AK��ߴ9�l�D�Wv�L4��-n@�.[�Ñ�%g:L)G^pK:M��]6Io�I;,��8nA[�\Р�dcL�#t5Y1
z���)����Բ�G����3�c��G3�����dqv ����B����kL�� ����}\�t�ŏ02ˠ�
糒�����wn�~Y4���.�� �	��'�:V�_�E���($Ivzx���b�����e���o�ُY�k�y�A[��=Z�h��o�+�mK	6�)͖Q ��F-�>��[�fw���.�;S|�G���~������!d0-*��`��Io�/�{"���^�CI@�ꞑ�����e�.����K;��U�l�������[��)��5�뛵x�1hͻ�c��6�h@�*�[��M�?�<LĮ_b1�빣�H��4�bG`�d�3v63=���A��ҧMha�1��7�KYs�U�� ���?�XB�-�8�[= 9���o�	 `�X��;~'����d?6�����<�+��qE�O|����c�,����^�L��ȅ\^��lQ��z��lG�ʟF�|�Û�J���I�W��3t���x1"��mh����@��^d��f>�Y�H�*RE���M�I��@�Iu�՘\�W0�)$L�-��2�&}�I�$��-l���o[�5���9iUO��=�T�#���<t�C�(����:����7 �LL���רW�!����@��m���r� �C�x,p�.IBԒ��%o�83��^�����b��͵a�Y�讽r���Xb�r�s D�xqL8o�X��<T�L�O�,U��������C��.����-�`vʮǸ2��Ӗ��!J���a k���E_u�P]`�g[R[�8��^�́=!f���x�\=j�m��l8��zu�	��s��aW�.R�����}~%D5���$��4i_<��~YzΘ�[���-�����t���1��[I�!�VD��c�j��yo��Y3��Hy���F��V�F�pB���g�%��"�_�Bї��)?������	S��m�=��
J$򍣸����D1�󥴔[�D5� ��x�ߧ���燿�+��h�a�ȶ����B�>�!�Ė�6*�Umd�|U5dH5�;@Z�hF��~���RE�7�8D4���n��l�(�P�s��ε+խ����ۮV#���wr�p�\QV�ZV��{��g9i�z�g��r�V���F.C
{.�
O�-3<��.ư~���6�d��l� ^m���4��A�A� �3Bd0o�K�|�9r��P�������������z3�}���WiT-��ӿ�X�=��{6�D�\�N�(�u"h�e8<=��a��i�N��?J[�诛ρrBQ����m��5D�I�3��I(z3,t�'�ʷ$�$����MG�9�0g�>D{/"�0��ľ;p�K�jo�=��h!� �4�o��-�E�I���Ymb^
�	`�L�G�������.7�w������L� �"���.�h���zfσ��	w3u�'��t��x1,2�ڎ�l���J�y�.���Ǝ�!��-Pp1v�$��\g��ԏN��5�?��t�n�H���_6SD�a�w������$���{~���jJ�7�KɌEP�Teރ}�%�A]���bR�LbG�
 =�h�<�������O��}nb��<v�{�V#�Pg|t��JG*�@���?Ц��>�f�b/�^�I�x�/?��#=��˰=ׅ�*�:��q�re�:�v�Z��k�P�<�!`��a����"�ʄ�EQ�"���)O �U��[�9�7��H[/���+J�B�zhW~d^�R��7igY�+~=>�XU O�E<C�AJ�U,�>�tSAt�bܜ�
��t��͎�׶A����eL���]�ae���l�����!���*�L�����csD3�&\���e>��p��Y.0��Mh�M���x�e�x�I���@�da�p��Kl�_�o�yZxq�� ���R"�\ͳ(>���Ǯ� v�vf����1��1������dd�ƨ�8?3&̅���� -���#���& ��x�`�}
r�����uA�@���7m2o�jJ�H誫d>sf�F#�%�Q�9H�Vҭ�ې0�E�w��$�c��˭āf½���p4]d3����?Vxa��aJ�C!����}���d���כ���%�dZ��ΰcQ��?���T%!���bRE�܏��a�1���~�x����bH@"a/*��	�\M]mBz���6h֧˼���V ����Zw%z:GM���C��>1���Z�,ث��X�9��oX���)�^e�P�u��O�t�!��?�S%^y��g�6�<��x�ۘ*�.4ˠ�����I��!7�IVE�}b}�{'��o'����.mh2��V��^}����f�!G��Ƒo8j�Y��~��⥳y�E]	���q��k :V��<�����*׀�v=)��}hN���E���놀􉤥��R��������E�P2��������Ǐ��T�9�`�~V�/] �X�]�w�Z
[fsuM��.my�.>h��2��Z=�v��q7a���ģ����W���S~�R�p'���I߆����ck<z�c�.�K���1z�\�p��r�{1���gWD������s����	2I���2헁}>nk��K��~�I9�&�fL���|s�xw˳�����Glމ�0�8�#xh�$"��_�	4)ɿ 1a8��#�l=&vK�B�F��8�`� ґ�d�tuN����0�W(�(H��gխ���b�����|�Đ`oʘ���c:1�A��m�Z��4l	rcY�'�b�Iﾥ�Pu�@H<h��@�8��B��*G����eэ�a�8���r�D���/�S?��	7�X9,L~"$UO$��}��rW&mx�XiTlBM�8��Ӌ���ȁ�<���!R�k��ca�����(m���i�~�])T�κ��YG����d!�T�Ȕm�4��؁��t��Q��m��U�m��ޒIZ9l�)���'s���ڬ�l*���Z���}rAƗ/�G��q�pUX�hf�{k���$*j�#�|_��	^�Y*:6�2��3��%��ɚy�a�l���[o��en^<���'��I�E�H�à���M�X2}���B���j��x�'��@�O���C�pȿ�&��<»N��j
�"��ޓc���r�8�y�J������l���A�_а�R�:��d�R�e?V���|�� Eq�Y�\���g��C;�Ɋ�a}'��C"�[?�I��G�����:�^0��}nE�5~����E�*Ť��g�e�uݷ�v
�ce�؃���#�P�k�ϧH��D���@ɥ	�|������=["��*C�����)�v!,e��%W����~��-db-�khkӀk��%[�&�R�&��E4�P�@�B�٠އ�5���sT���oD���+�_u��A,�|f�<8϶؂+�p�� {�&$�ʃ�	��	<�U�Kj����SC�:��(�"
@��-Y���?�5|+�?��v:�LeѮ�H�p�l�>���Y�㔡� �A����0a�X�K܁z�4+�c���.o����u�o����Y��a j���f�ꈻH��RX�Z�w�y�*�Ej��!����>[-DN��a���X3��|.�#*]%�pv��j<�z-,w�a�8��L
,����ٲ�8팧����-(�઎�H��o��5|�ٶ�=²�3<�qs,�/�-ͷ��͋E ��\k�#3�]R0W�9�"�x���b��ʣf%�
M��D���V��/������[�O�[�{Z�ǥ�Ա��ؚ���m�H��|�fd�}�XD����GI���J��*Y�e�����{WM��%�1����ۅ}8?�ek��`�TW5��e��u_?�V~ǚ-��2�U�������kY�*U1H a��p�� ,nk�4,=n�7
C�_�]R;�S� �h�TO	oz5�IZ����8;�V7{Y��Sq��稃����B��7�E��G���З�o���I5~�:Hx�S����y�<�X+�W��Z2"A e�5;P�4
�,5+TO��^�U%s��E|6��k��+��z�<��yI��
L��O���un�ϟ�&O�%a3B�K�!J�溛�E����%��P�9:���P3�_�h䏡���4�0�|�W[�O���ar+��7S�}������	�-,�bp��j�sd[)�Y��z/n� {�W��h�� >�j�@����~-*ۑ꟤��.���Un퓏�6�ѱ��^�|_�z�R
����w:Ѧ[9&S.mi�~��M�h�!*�h���-S�Ņ�g�3�B��������r����R��\HrB�-!�ݝ
�Vt��dc4��ٿ2CO��_�FT��i��Ʈ��7��Ǒ�n�L&���	��1'̥:?�7��`��Q�Wn@fG���8�_,����Pԋ�Ec}֠�?\�W���6� ^��V����sFЬ��m5lF�\����X38�.��zx➽`֐��A�����D��Q�w�ئ�u1����)�%���iaݗxuu���7Cx Ymѣ� ��'�>3�I[Y&N$<�
��EE�ًr�H>��4%�8�/7���ܟ�U��~Ì༷AIoh���̿�z~Q':�V�I��K�δ\*r����� �2�$��>f����"�ǅmxh���m����G�i39v��f��ƙ�!�$�

����ʸUA�з����k�(�7Z��?[�p2OW	��*W*(��5e�ÊKX#�k�=~a�x�~^L4R�E�B+ŭU ������]����>!~c*IA�>�Fs�L�R�+����+���o��||�U6ژ������ SFNS���^�/`�M����(�X2oԴ��W�,N�ՠ}��M��e�&���z�&�:6�T����L��v�I�?�L�� ���P}{�N���!��L�H�ݺ�PS��dH�^�[J�\9��ky�9lѪ3���Kw\�9�o����K�0�5��[����l&X��5q~I����W��I!র�Ca�3*��@�����?ů2.�/�N�N��~13�ԉO�:�8��ޙ,ی��k��:/�1�vw�k���$��qǄ0�{�'ͺGm-b�Qr��C1�dt,�R��wG�l�e���zNl�9���*���nȰ�{�!��Io�l��3��[֟���V2H�DL�/Y��M��s����"G�?긑�)X�>c�E�L�|n�[K{��b�����	�B�0��B>M��#���|_k�UR�3>�7 ����a������E��^�?������FK��dU}�+����08t��q�l��MÒ��H�y�r;'��9�_�{L�$}�0}T%��+0T��7	�0ڡ���5���6g|t���/�/5m�r�h|cl� к��ý���ym���+b�����A揌x���I�5�0>�����ܖ2"h��A�%+g=���z���P�M��{��#�B�(nL�Ⱦ3���z���U;佼��U�DȢ�O
�e;�t�K|�!������	-���T�c�)�5[��iX"\
�A�B'�Y��Xf���!�D�I���ٌt+ek��&z0�@%����o�qU��lR�`tG�)�U�"�u�����48�`kr{|Y%v���d���o�	��w��4z>��*}�k(������pݐ���)o�)�UC!?+(�nuc�7J�9�Y�ˀ�&>/,�=E�3��&���ɋ�^a���r�%�07X���U�M^��"u	Af!̤Atj]:7:�j�_6[.�0��u����n��&6>M?�*c��K���^X��Rse�ϔь�7C�ȝ���_�#�VX��0^,����
}[��?���������۪:�o�Gz���B�WH��`��!<>��j|���1,�g�5�tF���z��=f�#��6i9{��� ���{��ɞ~Ϧ�>���Y�����k��$��v����5��!h�wlH/2I����`�J�U����/��x��6�iѝ�Y3�H.W�&�D�߳x�˒��F����4�çc���Hx�e��3�7Ue�C�ZT�?K�h�ا��H#�**�,?��?�*�)v{#*��x���1�$�����Tk�\��5�痛y���Eum�P��g����jK.���?��	���یy��د�����q��oAN�9���}�fR���tJ|k�;�;4e�i��R\2�x�U�&����tiw��Ԍe����|�;����kKzq�>��x�\�_9�=
Ҟ� ��GR��������ɺ7���}���
���Vaʵ�K����`�.��k���v�2"x/���§x����,"�)��]���0� _{����ƈr�������DԎ�w�Lй넷Y �w'󛏞[��D�8I�ٱ�����`i=H@��.�ˣ�#��E��L���f�ј��\��L�Jeu���Q��9Q��"9��Ͳz+��њ�͛��>&���|_:���O!���VK;Gd>�� !.K ���yW�h�"s������9Q��F [�I�4C��ι�:�
�+�zG4dD<����̯4�Vy!�n�Rf��&�g��77P���{$�]�|u�P��rb�UX�WmR��%��[Q,���6��Ie0�f:�k�2���;Q6�Z�Q�<I$#��g���M_�R@�+�Ah�h_	��h�:����-*�ea�O�����{�E�����nܤA�Н��Y��k�G�GI��/�Q��]�K4����$�)�1��t�c�%�Xb��� a	�V�WbC���|oM�1��e��c]O
����u��`7ܙ�ni�L�����dL�Q���u#r�̍�օ���mApg��o�`���e���$�b�����=c�����Nln#�Aq�gD�U(�T���� ����d�L�ݭ<�M��}�"g���F1�K=���X��J{�u������|�=�n��C5x¸�+,y�(p�Ѓ�xD�+�9�Vx��)���Ĉ�; TnJ��#�C�X~�{��U>~C�5FN�2��i�\D�;)YY0��8��F��`mM�����L?ZFȻ�:��6hl� 	1��� ]�,�4x1��S�&�h|�u�p��Rdh7�X�ЎBX6G�핤��D��e$��5���GLU���;�����)��� ]�1\ޡC^��aqa��C�QB��,
�ٌ2�g~�B+��XA&�kZM�T���s�Im�?]��Q󝍪��K%��'j<'�h*��]vN��O���_P2O��Oڇ�%)�ٌc~���EEd�jN�l�Ѐ��`�cp����$W*�
.ӥ��f�6�7����׹�� ��LNDe}N���X����>-[d�ң�FbcǓt��[�[��X�*n��PS+uc���%F�r~�6JJ1� VP���֙����}^�TI��H7�qb���-��W��g�}e�h6r��U��Q�z����4�%،B�+<ݵN����x��=��Rx� �)��uV�.��P$E<h*|��C�,
����4��2i���a!Q��F��|.���Qm.��һx���ֆ��9�/���a��Q�7!�:2���E�}�{=���[B�
+��<�lΣ*��
;���t�2�3�e��|)b+T+�\���8�A}�a��>����qd��|i_��6�����(�^V�\F�k�6gr���E����S��q�2���b�A�<���5����aD#�V���k�5������T���nvN�z�$����P���e���̨	T�����Ѳ�Q!��7�hV�L�.��bE7;����ƜMݨ$�g[�%	&���%�	����p�;G'�-����n����MS�<�s��8���o�i�23}�<U���"Q�sd��\��.�� I1U,�޽%��`�5�f��{�r!ἁL���G�{$�q@ZE�1A�E+Һ����yŋ\�����SAm@�*x��K8�}���wl�T�!�#Z�Lb�����?�d��mM�K�gu{�T�ho� ��C�0<�#6�{�� ��8U͕X�(��$$��c�ع��dMD�.=���?�������5����rNA���U��a�VnxC�5d��Љ�;��Us�sÒ�� ��5Aˑ)����
)H\���F���U�|�ܤ��A��1ꮙ��ɴ�������0a�=h>��ծ�	8�t����b|rJ���B�����Ϊ̲Z��f�ZB?��Z%�m�Lq^�����IFe�X�W�b�{8p�\�׾t�J[i��8|�eI�%��.��쫍�P�h-�ՠM�m�~�塗�Fݵ�X����M�}q��.�jέ�!l��n��Z���EX� �_��)x7�������΋��4�P�?����d�Y~uPhENMR����&l�ML���pu�ٝG��GsJ���#��mM�ws��'k��U���!����F(�������,���>���
�1;�N��)����7ޱ���䇠)A�{KvU{<ħ�䓦 ֔轮�� ��'R%/w�!��h��4�((��w�.M�"0Nz�K��9�$��a�-�X�A�C�r�������87/iw��;]b� S(0QE͇nGK��h��1!s��5�M/=�͑�U�{5OӐ�;�Mt���F� ���G=���:�ܹ|���p��#Ye���E��2IT�w/�W���Z��E�� ?���ؘ�I*�3'�~�!)�ebc���Y������m:��8����s�/�>A�B���<���@�~��s <b��}bA��`��k���!���2������a��DH�sU���9Ř{ᬆ H$��	�uш�ZS�J��Ro�Qݣgb�=�Eu�>��� �k�Դz��$2F�(�?68�r�U��~�WZ���j�X	���`�%WZ�'%:��:��B�d���t���]�g�w�i�\�_t�<j�ǐѳd��`���V����B2���:�3�Q�K��Y���Ś�.wf3.򴙐���c��w�����V��{�0?�k���֪%Y�8s֥�DO��?�me<*h5��hLN[���9a֌ @��NL�����.�؈��:a�|*�?,����=��횃#�Uv���_�C��,�L5����ٮ|���r(�m�V�2��SK�0��Ax�sɻ�0n��w����HZ8����ՀH��Mz�-�J�������czE�8s��l0i�߲~�����yª>H�H)��D|%������?�4��#�_>Dyrr��m��I����]9M�|����o��u&O8�o�}��M8�g��,M�i��]��H?*F<�gD[�|���S�j�`oX���͟h�g�g�$�:�2p$@u����ӵ
����q9��W���T��x��ʄ @�F4sN	շc>m�wt��Ű�C��j��=mʶ��"��Ĝ��K���,��^�q�x�3���X&�p��/�8�����\�5םEkBsH;�pѰ	y3q7r��/2��`3��l
�F{�X�X<���o��=�z��Y�c�*F�z8e}������j�j�Hd�cTU\Ns��H�	Obw���p#Q�}@����8�lv�?^;��vO2@�M	�7�L��:��v��_��6����Z�W?P��% ��?z��u����+��"��囧ژ-�R9<���������~��Ɇh���(<d��@�^��`��Q;��*���:M��98�w�/ƃe�u�)���A�ü;1�0�<���`���`P����w�2��<D΍�� i6�]�NP�Ҡ�i�A����:�]�B;�4oq[�W�������$��y���pK���v�|���������p_+���IK�&;�"�E�Ɍ��^��b�U[:��¾H@��mxp� e�&�W���TJ���������z@^$L�*�ɦ�rkEW���9Sa�U������62j+۲w5�BHZ&1I���rîE
y�=�=��_�(��OC'W���v���ˠ���E�������
�N8p;�vG	�ٻո%�S����X"�Ɗ���`�rt]��R���Ҝ�b�9U��5����rN�͕ba
A�{'����&��;��F����/aɗ�7~��L�W�K����j	����ۣ�ɤ�8d&�
a����ع����G���:|@Y0�?='��^{�G��xc�6�,I3�==qY
#�N:��n~�;��ن��59��g�b;u��A]$����k�稘q<xI9����6�t�蓁�\����g �T��'��3��8�����s�^iJ�M��{4rNw��*��A�m�z$�u�u��w���^Xm�eS����?J嘇58e���e?W��н��7�i��f��a;�Ǔu��O���f�M:��Q��H�o�|$�1Q�3m�2w�g�&��vm��b*d��5m�.��a��
^�٦7�F�ޱ�Oϓ8�;��{7�����z���)�e���*Q����(�y��?LʕW��!�2�a+Ó�k�o�/�r(��!d��m�8��8��,�>��O�PM��X�;��R��N~�[k�Qx�m1cG��w��a�4�:�O�����6Ǯ���N%s�Pti�m�����ŲS�>��n�����ػn\�Q���� ��ԍT���;Pc<F_�BpU��������coA��Z c�^�#�c���{��u?)�uZO��g�6����~�%�~Ov� ��_`�Є��y�/S;�`sB�"��ç�������*�:�Ff�3�+�C�Z�!��ّ�4G|�S�@"龱� x�O� t-a��-˛~b$</�]`tI�W?�ڏ��%-zb�]��* 8��(����芏߽�a�}{qC�N�b�,5�j]���B =Hw3���e���3��LVS��Q�"C��5uw̳�@����Q4q�����8~r�4�
��>�G@�4Q�y�C�Q9|>N��_��)����T�����F�mj8��d�&rq>�C��w��Y#ؽ'.��1x�9x��Й�8�#���DcJ;n2S�6��W�2#�7��������f	���A6X�����uB#��K`J�_�9m���5�tOzf�r�.BO�i~~��4@c%_r�x�����'��G��	�f��5��<$N�Q��N��@�����S!��P�7K��CT��y �L7����>�*xu�w�T�:USK�����]�%���ri"�C��EgG���h`���3p��Z*�v���Nr�Eb]a�uF��Z�eN�B�}7�&Y^F{�����wwP_p5��UCRf�����)���H=��s�z�_MS �'B��$����X������th��/=�]�_8;��4�NT�V\%��;fY�j�i�c�j�#�=�,<�@�7 ���� }w'$��Tx��E*ҁ/_��E�s.�<>�\0�~��x8Jy�:l������Fj�L�c+�_��vn��;�̚�i�7mZ��Yٺ��h�Ac�N���y�$��j(n9�Ѕ���?�m�i��L�~��{&�|a�0?M$�v_�8��*�
;�[��(�v[�ɖrz{Z��3�Ap���=k�����Z[72e0��`���I�6�2�i`1~Q��Ϊ�3U�+�r�,&�8��`�M��Y�������>D%�F��\c� O)��;�`�Z���RNKk��[gD��N�^
T+Rm��r�rhC@�����{���^!]�ϯq0Y��,�qMU��\�����=�˳Ԍ�g�����C�gYO��@`-ho�OI�<pBGaj'�l�b9Z����bu�]m�YV4��Ҳy�SYܞ]�N�%���`���}�@^俙p��!�5c�1G`JyEn��;)OI,"� ksN9I����:�*ts_[	�����2�Շ�\����f?;c��I�;Jn��e[)���$�B'26h�4յ���B��_�~�SV���u>�2[7� ��9z��z���C��R(��[X�r���*)��kyt�ľS�ڟ
�{��Ƥ�Y_S�@=׼rK-���-TUs�Ǔ)�a>B�6�n��u�~��Sf.�A�Sqy=�q�G��+��p��d��_zB������(�3?�Խ��l�Y�Q���/*�g�<vg	��D,�n�Kۘl|�/�t�i 6N1�h�QWL�x�%f2�IŃN�z�^�F��l��[�F�H�p�Gr���@�!v�t�_�e�_]�sO�0X?F#�$N��3䡯���'ͺޱ-�@9x}���L���h���� �p���*���	���7�A�����������TϜpwvJ�ВE�:����1��;g��Wm�x^�#�AC�nnh�^fz�'gi�4�'�!�ڭ7jfy+��Q~{�.�`@���Ū�Q���U!���-��qT��RE♉�y�x������D����,k�'����6��kt���6�l5��gy[����˔�Ia�Ͳ,�ąT���px��_�"H�h�2]��4^�|Lk"UH�A�<���oQjsh�W&k�T�,䤅-	B\\h_4�iy1G5c���,,���74L
��k��R��� �A3�Xf���B�b?n;���ȶ�\ ���#xu8�T�`1��M�}^�^��vΰs�i4u=7Lh�1�����ǂed1s�Z�>�]r����Y�i�m��b,�hb�r�z�a�(D��E���d��q
��dD~��vIc|�ڡ�SaC��D��a�^%�N�C(}��ǚwq���\��*�]7��1Mt�=�j�S���Tj�Bv=���o�Ηt�`g���V����\�b/N�D/�������p^P�v�'�՘�]<h=��䇖S.53V��Q.��U�l}Y�9�rh�~�iZD3k( �|S8��YV�P�gۘ��ja�A����E�B4��p��ɛ�]/�k��Z!�F���ւ-��������y6,.	�׿���S<�u���;"�<|���3í�7ʤ·H��At��MY�����u)e"r�VU��B}$cǐ5����ˋwV`C�*<v��姥����ZV^��Ù��j{$�ty�`&�'�UyB����Y���I��,��@�hq�[!���J��ew���],���!a��s���B<��%3Εǋ�Sp �L5n~^�Г���v����lX}o�\�:�h�>޾̨Y�g#t
X��A��qKf�X���*���F��sȌpk��(��6bp�ݭ�HT��Ta����/��s�D~��6�}U�Oh.M�U	�f�hP�C�?���{Ɍ�O[��X����W�3�\̰�A�J>+�r��@��r�n;�����{�U�Z���x����Ѣ�ǣ�K��
=�i���/����/�^�])0�軜M_!���������M�9�iR�R;X�K��Wd}7��.�	�L��(��y@G��u/؁C�Pߊ���D��S�:`;��O�-�ה�ūeղ�_�U����~�n��u�=�@_[�"V��wv^��0�nX��?�9����#��x����w�Hn~8���²+�x/��lZZϱ F�T-��_������ˊ�|��=��BܙT��+D q�������r��V�`(�U��4�p��k/A�m�4	E�5�Q��Ԧ�A�8�ʅ�i�ۈa��x�Pm2d\�=�;��ӭ2��,hj�2�E�F��/Ό�?���,
|�/��@����0Ӭۆ���imKXr��Ma[�8x���p���W-L��<q�;�ǔ�*�$�޿���e/���lHn����>�1��z�1�2����靂\� �L\����a����m�/-!��H˔�u�@$v�e��]�
��	P�_�
dg�b���<R�T�̣[v�	M_�$�\����"!�wws�,�{�x�d�˳#�_h�w�&Q��ź�ՕhY���3@^kF�@����|���d!6W!��B��`�nbQ̣>�<��e���ǰ�*�^��g�e���֣Lb"ui�
�:~��-FC��䠝V��qT�D?��9 ��s�����<o@�!(h{��ETN:�5�����h��� �l����'��ɛ8`ҭ����Ea�t[ɑ���~�:O�e 9ܷL:�9��<���:SK�X�{�GaG�d�}�z�u�Ի��R3�B�9�ɻG[��p��c�&T�Y�Y�1�Lz��h��I�Z�7ڼ�Rr���s���	"���>o���A�a��9T�Lk$Jh�����n�ﶕ T��x_<0��G,n���e%��-E���mSߴbmY��p�'�$��Հ��A��;�jsF!g�"+PY����
�	
?����/^�q���V���P�����~xrq���%��G<�?]�#� #��l^ωJ�R�_��sM��ݩ/����k����a5���t���V�NQ a�J�3�d`�n��ԍ��2��GisG}K15��)�Y�Xh�Pp� �$C�����8�.����gzӢg���[Ʃ���z�R؂`ia�C��S���[��?S3��┲�'�6A��������,z���2��Y��ea]aJ��
��)�̾?.�fR�+n3��f�vA�7��q��*���o#p�U�F\���R��H^>�KN���X�&�p�&���߻����'���� ^���P�����K��Q�1vң:B\x~r��%�ՎX�f>��-�Ӗ���T:��S����~b��5������o���i:�ǩ��a#q{2��u;��g/P)�#ر�hqm�������ZA	��r˜�w��`�6&�M���m1���h��ֲ2,��T����c8N�/��6��̧5H�I�h�� �E_����]s�V��&�	��'!��B�'������G(XX~�dAoT��7���[�%?���y��Z?�|��q�M2r��H���h�)P��/����NĘ��nPt��HS�0�d�
�Y�p�LJ�řK��~�o����A<h���x��="=י����p0��v�6"6r�'h�lܡ�� ��K(\��wm{�'y�f��8Pnq�_���%ac�cp_+>ō��≞�T�\�Qe]s	Ns�E�Q�M� �8tpqk��j�)���E �h�ٹ�R��d�nP�� ��5}>G�~N9�؏�~Y��w02t��McO�3̍���T�vqqz ���m�`�5���\\��{�a)Ә�@D8����Z��ᬊ`Sop;�.�r�qY궏�^��Q�9��~z�p�. ���Q�-r��0�����GҼ������@y�|��gd_��;�PK�����W����(ޕ�yEl�b�T�' �Wo.N�ӉCo���+s�x;]�(���F�R�4�^5|V��|L��-k�����qrz+*+��C0vʋhЬn;W$$$sj"�/��@��!��Lc4�<I�������Nx�\�6����n��V��d��������P!�qmwW�*�O2ex<I!������sv���RFE/5� v|�̟[X�D;Kg�}�ڦ�� �Q���v���Æ��+j�M�ρI�"T1�W���Oy��C�v	N�����*���BѢL���˴����
�Y@#*�릗0�e
�6��Q�J�<fP���4��	�ޛ�Y:��'"�J��3�t�Wy�z����g%{�[��ý�3貈�u�It�3���t�Ǹͬ�Ĥ��g�N�斱�. ���*�{Rɒھ�i��E�d^���X���֖�����E����u�d��9F����Ȃ��T��S== W���l��;��	ͱ�/��/���v��1!�>u�P.�fB�zc@��y��5w��;"O0��%�kU�dB��sX�z��ps0sC@���W�8Y�Z��!�}�mZ�,�mK�:���%H&��� t��ԕ�5���8��IeDg��56�n������* ��nc�07���}__�Л~ŋ��q�.�+p=o��������d�Ь��'���
hh���E����U	ꎇK�!�����g�	�NK�>ɔF;���TiK_�t�;��H�c�
Q��>H�a�b8��yx��׭'X��̽����Ȑ�׺��BS��p��������8�}3H�+�����ˀT��^�=oÜxƈ���)�9$]�tI�H"<%Mp�����ȗ�'1�]��.6��d���)��g+��#ơ� kv��w�pcx���28c���qWu��l�-�R�n��]���{������1�h�o@ZXsI�`Ś�B��B#�lsg?�b����G�y!o�o��(�n�����\����/ �V�#���Yr���n������El��7����_Ok'ѯ�$�x�-X+�{ �6s�B�z��NY��9�oc���ȘmU��S��q��}��#:|*�Ū�6�cl�$?]1������eq�h؛+r�d�=�6?�/\������{��>�q0��2r`i�$��$?��ى�(R�E9��-��?��T�n�y�Qs{T�����W��О=�{o7����4��g�H�e��*�'�(&�oY3�f��s�}�>�`U��G�/�|�1��P�f�mj&VY^?Hk�Y��j��_��(^J%qk��4�="U��0�(���g�g����H?jq�Аb>GK��V�]Xn����K�(2�8X_���c��E�ra�G59J�~S3ј�]��`L����5�Q�����j��9���E�8������[�R�a�&ﶌ��t�~ǜB9�`�������B��0�86&�����4�.��>�/I�B~%̧��V����ԭ���v�)�G�~��o�M+��VV�
s��`�����6˕^�~~����sT��iN����+��� ]�?m9�n"iV[����Я_s� q�Z��0��:g��edB��՜�]�퓡���ؽ��Ҫ��-ǽ��Ɛ�F�'�xU�6	��
.;�,2��I����(3���}c��1n�2-���ʀ� 0�Q��ؼj�"w��ك��!p��Ҕ-Z�A������Yh���B&$����0���=OҐp�zc��0%���~��y�˪����E������)�9P��c���O(S�\��!��3�&�X=��mA��tڃ�'��*(�b��A�R#���#��5
 ��q�i�@eXMC��x�#�w������fp��!���+�U+�p�km�8��*�s�}�$sM ��/��A=[�heu�1�;ԫ�𢌗"����[6�Q�"\ h@���
�!��tɏ\���.4����!D�*�v�Ŀ�nL��iC���YYe�1g��~�A����E�ƞ�ſI6����`����t��F��8�$N�ꎩ��F���:Ǧ�Pl�C~㈴nx��	�j.L�.��H���Њ��z���}��� ��*�r~�
��6�L2d,��[o�J�j)Pao{w��z�r8A3���*N���[���j��&��>w_&іތ�p���A��5��W^(ɘ��9ڠ�adg�!sXZ�.��V�44ܸ��i��O���`C�M�{B��9/�x�5h���W%J����Ϳ�O��{��T�MB7��.�������"�����L�91Qٿy�vGPd*b�)��>nS�X�R.�ϧ�:� v������ͨZB�I2��<��ק�t|)���	vL�h��A�)y�ń�{lA5���u��-��^�S>{�*�x�Lۓd�y�������(ƈ������JU�j}=ṝ�9J��卻��R�ȕ�lT���ɱ�*"$���>�}i����fp��Q�mV�s:�[WF\p6�O-1����$������	x�dGj�SI!NP)ޟ������j2����՛~��h��s�-�^d7�pnjmb��͘za	ƾ�}r�f��� -ᝆ���[�e�����o�Qz�6�4ob��Jr<�/pc�嬠��=��jb��Nܧ:�{�~��n6�l���J�5�F��z����-��ZޫP���i�&w9���%�Q�s( Fr���vrs[M�H�=sW�6jOг��nX���ɼ\/��?��.?�P+,ϧ{p�x�)ȱ�VfЪ�Iu
�y��W#}�N�"*n�T��+,Jg8&�Ǭ%ǡ�V[��A?��U�f.h�dƎQ�#����D\b9T����;J،{-@���W�+%"��_sb9QA�`>\I�<�)#�]�����o8_�-�iu=^��T�y��-�+��BV��.��벥d4��x��R�f`��i }�����_a���b�)�w�����a/9i�/��z��REK�h�F(���@8;q���<ve�Ȏ�FD�����|vRZJ��a�O��(�Z�l�{i�.�0��Z{!���e�S�ssq?si���3�դ���G3���0�}F�C4�)]�:���)!�J�|�i���rzNҙ�A�AB�ǈ{;��@�O�KpH�9�V3�@�h�G���N`�FS]׏r���\�| ��M�jW�.]P��G�R�����*�;k�E+7���l�V���,��q�D�r��A/�'������r�<6��`�R
��(������&b�3l��/�ΟeEV
����z-�ُJ�PnBF0��8�u �����;�H��U9�vgD8����mO.�c�k���ʰE�M)M=?;E��$�p�m�8lg�3��NП?��׊��� ��Lt[s۹g"��ʌD�`�ș�lVBK�:O�&���J�(q�(�YrH���Y����K͈�e?����軰�.~0�P�$��BJ��I�#|],`@�[Y�T�RO���㎌X�{r���Z��[~�"����ݓ��z�\�]��-����֭���(���a�S�N����4����V��}U�m��a%��qh滢�R��Bϴ�]����9&Joa] ��|%�����v���ʲN��m8xp�!�x��b#��VU)ʴl�G�2SmY�z�  A��R�61w��>v)��c�k��G��U�d	!�u;%M�2O4]��t+���L���<t�׶��gli������p9|ps�n�(�ń��R��XD��
_&Z2c��Za�=f�/!�[��I�yȡ?�_�+��n�Ȟ�f�fQ��p�ӯ�\~F���5K�j����t� �Ghۀ�L�D��xLT	#e�����a%�Ld��Y��f=�v{�"����C�1b&�=�)���XGU->�H�A���?�y��p�yWpy�9��]
�y��]>��Oh!�V#�dtu�����yj<�y�u�^m�OYڣn|�pQn9��r�C��z�z��Z�L�Ɔd���:���|��P�	^Dq�Lz�ik��	o��\�ç^{Y%.r<��tM�5]~�S*yL�MTR8��o��%X��Q�t�����xE4����$�Xm��-�4��h(�s����9k��~.s�L�d�3�la,��"��������ˍ6?���a����bi�Y8�n�B#?z:4D��1��tg�^౛���2����"dwA�!ף��93�S�����j?���FJ�����U"�����������
���D��!�aM�p�U���h�,�O����(@x�Xϸ'�� SaX_5����7�6$�F����L	p[�g�l �G��M}��ْ�%!���@خ��-^]*�|n+���_�LK�:<V��u�!hն�M����
��9�����7�8;~"�//�)��I�W�8��Dt옯�I]pJ�]Ղ����F�	`�{~�	P��}���Sh:d˒�?!�?�Dc��dA���Q���T�`�<X� ��ѹ-m���:4��@r��B�yVsB�<[�0�7 �[�h�+�D�g�fw��O�/C�[s�B��-�-���3݊�c{�}!65S��F��db]��R4:��be�w	=�=�p`1�?�j�@�oM"q�f.�?�j�5K�l�(��7Ĭ2���|\:DTT��'v��9����!Ui�����ק'�LS�"�5gy}�Ķ�q��!u�뿠C �k��m��t�:�~��DQ5�\�)�"~�pÇ�w��N�q@'�����ؒ�䤑�t� �NС�\?�=��t�[�=>J����u��~C K��M{/�	��1#��?c�#�˕e9�f���X6{߲DظL�4p_�	�Z�����&7y�[�eᴂ��$$B�sq���|k���:�	���+J��%�X�L^2���'՝�;�t�hp�u���X�Ћ�֗{  g�+�E+�#�cp��m? %�<m�s�
���%��_vF"7�:��;:������Si
x>{1�1��#��������]��^h�ݟK;��?"
o��4d�t���,=z;�G�#��v����U�*��%K�9X�s��+Gƿ9Lw ~^��S�Va`'l��[t�o����x�&W���&�(���S-45�s;h֘_�Δ�#��˞O+�-�����D�d���"؏!���T����Nz����D�B4�`�D���UW/��8�L;Qq8���+�ҺF���&���U$ʕ\.�@%���@^��y+��1���55��|�u��U��&�HX*K�V�|�T'6F�����f���%�>�����V0:�������e����K"2�)l���|r�,ٸ
�+r�G����h�ߣ8�#�0�т��}{\�(�  qi��yZ��%�'˘�x�u=~Wp:[r��@���� 1���;�4B�|� �h��;>�����m��v�J�OöIPH������~Dv�_��&�T:��M"l��� {8*�-{�<�B��L��*�{fAYzwW�/5)�­UX.Z�f/R�E���DT�u9���_��jPϕ�������K���p���Y��8ߌ�Q6Ǧ�-]I�S�ME1�QU]�@�4��e������ƕ�ӌG~���;X$��-[=�'}��Q]$�m����C�/2Y6�F�7Di����׌���U����OZ���<��퐬�^����>�7%� �Lu[t�Hlt���*�D�ͱU��Epݰ�Rȁ~������D�Oc�`Ϻ.h��|;�w/F��<�0��I.)e1w47>:�Z�=�yY�3�9�HD.��p���=A�3+\�,j��Y�� ��U���Y� �hk�����E�3_�A��q��m�,�MFI����֠fz�g�V�G\]�_V<����"qX��Ȣ*yTk�B(�%Yߏ_8�GVc 2&W�c:�6����2��G񬫾ڽ6hQ_^V5d��A�tV��_|:N�=���C,������1�뷙=��VT�
�L[/W��G�����v����,�nL�D��A��v���Rq�N�y"uG�I��#�ۨp�[|���%����g~#�����^�
f����|.�O�qV	�m��+wن� n�ÜE���A�k�5B�%Ms^���X�G^"���3�Q�	�wi�_����x���x��%3�����CN���/�*ćyě?�ԟ]�eG�W� �wH�g��RR9%	(m0������=Tf,�7�q���ܠ�#6Rh��C���׊��Y��h��t��~H��_Q���o���ϥ�O�f�Ű��Lj��R�s��^	�ϗ�PY�B!���A��rw6$�Ek�ϸ��� �����β��Ug�J��8���b�vDv�~ t%��Xm���Nh�w��5�����6��%��3���WDMҀ �:�u�!�z����i�ӹ�:%F�˖��TaR�4�����=w~���pT��G�$���R��G����'`gH��� 5~���}7m��r8�ɞc
��N�����P;�OZn���[�b�z{���x�xY���J�F��A.@|���UBp�Cb���A
�*�%�g���c��|��O�Z�1�Ȇ[+@�XƓ�`{���/��:H�;� u^ĝV'+�nN�#�y�����zc�yc�� -�f~��iu�M�O��ϊ��+q}�몭�����'4LPca�0�����K����!u�~��C�o"��㵒�N���F$�򧞨���߂h���3��s�:���'1�9��R"XqV�wWS:��!XzQ�= rێq�^��^�8�%M�����OAv��ǖ��")�]�N�ݑ��|����v�P	6������A�y2D�h��H'?�R�NT�HF�Z���z��]�J��Aw�����l��AX�d�4D����xB���������ބ�Vk���R�yK���+h@� ǩ����X9�`S5���,�7��>�(8e��ғxϛ���gy� �&���w�I�X���gM��I��O��!�(h�76V7��)u��`��]�n��Ƅ̓��3U��nř3-�[N=��)�P*��M��o:ō4��J�`� hh6p�ֿ���+��yKB��:|�Fd�i��eE�2�/m��Z<��A�a�k4�U�%�}^Q$�Ac��������:�gQ˯:�Q�qx��I���E����F��R&�&ii;��(ӱV|���Li֓rV��#������+�[-�4ʴ;���:�w�"��o�J�yzb��q����61��?na��}��]BwG�TM^�T3��fc�O����:\\�K�}s -�ʫ�MC��9�
���I"��(/X�X�D���B�g���p̀�Ho���˽Sq�G�E�9�7�C�A��Թ�y��H�:˵6�I`��͐��z����#
���g�1/k,>�h�SB3Ю{�ϴ&R��HH�? ���� M����܁�����(�T���\O��d
����(��d ��iE3�	&xP�s�H~��Y�Ƿ�w�)DH!"%&ujY ����|R� ���w���"��&�P����/�ᧅ�[����i�7A��;��I���O̾��]��ߢ��L��{��D�C��A�6�H�Y���M�6Q��2���@�@ע	C�S�kI|���ޜ���	-cL���x����`Տ�u��#y���V�^���f��)��S��	T�\Ҩ(S�y�huӷI�9v�+��EN_���{Z�.|V����_�.�%�v��|��p?Ҷ���{jX����x@�l�  �e%щ��K�ޘ�����|�:�[%pW~�z4kEEd����`ze4k���֔�Jo�������>3����o<�d�v�8��,ʅ.ݦ��&p7M/��\2�ZH�N���A�>�a�x�%b'��� llXGZ���-֪�m�Ps��ƴ*�Qw�b#�E���T$��z]�0MuV�-L��y�i���`�3ᙲe-�bG����m�Z�9T�귕�@����g�<���^}N�?��0G�c�fhkp0/�����|��E�����A*_���,�'�
�ŵv���r NH��D\�s�"c�IJ@D�퀒��������=h����q�L��'�޴.�1�43v��of/�M���a��P�Ӥ�k%3x_	Ps+���ہ�[K�3��ܔrg�p }W��և�'����ń��Gi9�	�qa�	m楊(�:��������EK4�a�+;��X�U&)ڏKt> ��s���M	�(��T���P�l����M*��e�F�;��I9��$�+K���!���%맱E�0�mo`�B=$>P��KdV&Nf43˄O�9E͘�Ǫ�Y�N�="����!�].����]�#�þ�"�_�q_��z4C�ۘ&��'S�� ��3���ld��,`���z;�ߵ�̬y>�R�me�5�E�Y�+�K��r�	��m�S�����ȧ��&�fR��[�
�uL�&B��̢�	�\THm|d�}r�YJ!��E�7���ğ|���f <3j���+��ު&V0f�"6*+vu���_V��u�T�R��ɧ:Of�zC+"��;vV)I%���d�$6�^�V"�����Accݬ%	*�^a�c��,y��`�Ĉ�k�A�kc#�:;`?�d���ݯ���Н�ُsL�F�ou�.ݜ���=�SS~�������5�tB����P�c�T��9�J7�Pw���XB�<d3��xu���8��j��[v<Ӝބ�����=��X���֊��	-�X��:ug�2������(��|E�GSp�>�G@`����P��y�=����4���L*�!�Y�؅�{�C7<O�q�H-tR��_���i����!2����=�Aa��~_��!P�w0#�F�����.:�h`�U 0�����Ǻq������F20g�߉@�����}�y��SO���@֓f+��g��8H�R�S��Z⹯�����{�O�j\����-T��0��Ɇ��H�t1�?>�,���l���w�ܘ�������紵��۞e������:m�nupAb�����jB�JA[������(̞T�gߘ>��h'S���L)v��;�?���![�EI8���)���J8��1T"��.?vm�uA̚U�j�����UQٸ�+�o��D�IQ'�� 9V{s�f?�'NJt����9�"��~�x�
��h�awE�]	���n�(���C��G�zMr~~v:R�<��9�v�MێT�5��3�O��*�����v��6G��q5;�����D$�i����ڋ�p:U-3��+v���#DsB�H(	�3��/�1)n�2��:�m=��M��<�Xj���M�?K�U�G�H���a��G#�I'����dJxTwU���,�!�Jh-o3`=��T�����I��P�͓)�r��S�sx_��3��֕/�	E����Wt��&�Ϭ�Lq5�d��ٜ^_Ag�S0�$��A�����V!��l�6�t]Hh�9u>���Afh;���"cl ��TSϤ�x_2۾�m3� >�p���,�tJ���M�bsk�C,i��cc褑�|{����Y7��WW^��e��
C'��t/2M}F��U7��~JȈw%rǶW�~d���g����V�3�Q���Kih�n�-���ɿ�������ۭ�g��cNoT�w���1�~l��(�8�B�qG3��x��&��?���h��
�	���[�#��K'��L� ]DR���~>�$;r�!��=/UT��J�v�5�Sb���n���l�(I�}�#Y8Ea�P��	��ik	�,Z�)�Q���f��6��:Ro�Gۊ�p`�0;�صU��oaԧ(�{e��=������yC�D��=��{��z�<�u35�0�fnw0a�M�s�ܳ�$Z��Azz��Q��+���g�����9d�+
Ȣ�Sk��|�-�!�`ӡ6�y�����Dt��*O��h�z���\�هJ�Yv`�����C�p�.���"YF�9�^�\,��{�"��6˿���|
�+a�|�e�H�v�f����tܥe5�y�(�{�#��([��� ^>��6?u�^��~�1�w�H���Ʌ����7�B(uU���(�5�%�֏���Y�O��*�[�Kw��KUŜ��\x��!2ڳ�C��*�V3�[[����?
���K8:1d���t����֦W����?���o
,��z��I����� ��I���(t	�*�@Y1�$�-ox!��~�������~&ι2�5���B����* ��N���vB1��a@Ml������ ��0�'�{GFg�4���Zf�"]g:Rlt�ڒ,�i>	��9A�,����#|�J�Ǧȿ�xEг��/^\�)e՜�2�*�3a���#�2��s���R�;=�n]���(�>BUGi��my�f#���l;���"�i�����hp�ܐ'�0X�nη��z���@ꎝ|��@ś�Z�8"��)9��pF�b����L���Х��Qt��&�^&n�&!#4�3_��ηr��ba䗣d'(g~ܫ[	9�^V��-J&��w��τ�앿���e�TO�Oa�[�oх�b�����kZ�8���?;�#-�b�X�w��o�^%4ܳ�Gq���A� Aq�Møܽ�v����_h�?�����Cبz����!:���V�U﬑���q�g(�&� ���lV;�L�Z'�G����s�l���ٿ��E͌����T5�M�.�I�I���ĺ���m���F�.ѧ��`A��.�*��_tJ~c+^~ۂ�,S/�oպ�2���-�<��ה�1�� 5q�Ǖ�V�-Fe����1��
��"��ͥYw�L_�v�-y�0��О�}�3�t s���3�D|=�f�~�TF�8��V�yc"�T[��_�|�����}]� �'q�L�_� g�u��5&�"�-k	;���-�����mKV�i�}��!"��^�WP�(�'8�OF͆J���.�؂v���f���"�;T/�B��)a0�,!|_[��άA�ax�'��W0�|Bt�$�F ������V;�P��|�~tѽɜ��;����x<l>��W����n(A�4�Ky����t���!�@�9�$���'�H$2��ޯ�R����5�)PV���H�a�h&�R�;3�����[�U+E����g�g%'Ծ��E�bB�����vֺ&��-�s ӓ���DX����D%�P-:�Y�3���׫~7���eM>�E3��
�&��T�s��g�y�ڳ9x{m��I��K����zɢ	���l%�+����X	��Q>$��U6���k�{�-O�Lr�@�jӗ��(EǷ`N��f�d�W�=gYW�	�r������4�P�~paNZNTE
�-���&�q	,�k)j�>"x�&�	fzHmC�$���c�����1H'��qk'�a>�#-��jq��Cl�b�\g������/e<bSr;P���; '��|�b
�6[�<��G����!D�P���H��`�U�=Oә\��������Uۅ��_����++,�k�!�T̃��/��n]$�)}yDn����m����glr�R{�{�@>�Y͇'����:��Z���9K����� 
ь�:�1QB���䴣�j��l*m���v@�[�rg�I���������_�"��c�>	��׷:B�4�	*Lw`)x=�M'e�̓z�~�8�w�q���*j9��ua]@���!�>�ޥh�������OI�o��`-���a���3�1�w���0.��sr~t�?&���݂ð�߮�>"�Vл�~�Q> �?�nY�ݫ!g�����N蹄�s(R2�Jsm]f�Hp�Y�^@{������82oEm��T�Ie���S��-5����GN�1�+��a��Q$� ��o���(�����~Ϲ:ݐJttsRx����G|ɼX	nN�-��U����H����Ju�<pS )�҅��SpZӝ�=a_а�+9�t�n��;g.��n\�7��!@�`a%���N0+�1s�51��<�&��3�L�ys�L,��eH��~�vp��Q��G���RtY��J����GVuG�-�'�V��_I�e<�( dLR�̒�����?l�z�xK��� �Y~4_�;v� �^W�z�V�.�=���k e"Z�TȠ3T2ī�ψ-�.�Zu�0e�Q<�H����#Az�PZR���e8���2=_n�	����:�5k=i[]��D�M%��P@�J3���SӞ@���)�:���(3կƺ�E{�3FF�G<��m���#�vk���B�k�`J�ַ3���?;O�?�hv�@�<��C�{�!|ׁIޫ�+F��B]��m���rF�5��	�*�>��Eb�̒'���̈́V��z&ա�4�?��f�Lcx�`�@�!�|$�/���ê˙��+z$��_]53lW��S��Mrv��Gj���I�B�i#~�Zi
���[����)���W�D�� �[&�.����U�,���0�7Ċ�K}�k5�k9�� �U��҉�t�t���Y�{�� ��ĬM:iz^�����y��w������[l�f�]q�?�+Ux���mθF�՝浛 /��Ӑ�!��W �����8�$����3*=���6���LC�O����m��Bh�X�'�{CF�V>���w���Җ�F�9SLF�B2)��E�њn�ԓ�<������<��-�7*Y�]<my��D.�(e�n�e_g�����|9}u���WSd������)R�/�$Pn�ϘZ� :#a��\�I�� �<0�$@,��o�Y��T?�L���X����V���̄��∯��^o���/B�E-/}w���uO����z;�&�ܬ�f'y��	��ci��Z�7���F��������3s�~�XD�� ��6��Z��m�;���Btbņ|����OF��� ?�\sE����'�F�!D9%W�3�$֛�Q�̶���t��"�����rh��h+���+)�J�%� ���؅�
��S�A�x4q]�¯�k�vCE-�X<{'����l��oz������FA������$>�+�Qb�(��E��,-vL�l�����\J(k�N��b�W��^�C��Oշi��:`�7���?�r8� 8n��3#�w�Xo��#�%�Fo��$� U��'���T���~��O@��b���<�6���tXy.�j�7��W�Q�����,/p9��T�\֫�0ϸ2*���6�B��^�c1,��6�c֙{ڤ��+hiIuL�X�~�Iy��!Ĳ*OY��Y����Br�sk�� �<��(Z�x�X�\��׎�����&K}=��`T/i�v�,gB�\n���q�0�^����p���h��z�m/;�\V����zhN(�!��9�����M���ѷ�n�Hܱ�A�l��8%�_���@�1��经@�)�.��|�R&ߥ� xH/5�����!��l��1��9�4��V���#�7���RRћ;���zee�K��=
�
��2�:�^\�6zI5yI  gy�Ef5���/B��at�iBCx[-�ۻ6��}�� ��O,q�{���@� 4^���[;�G/zdY'����l��_w�o�F��%U4�/����EO����J4���b��B{� ^�n1N��G� �p{��0<3k#��d�'td��t�4*����q����P �v���=��
�_Vx�ui�G8��k�K���>Kq	����L�S���wFu�d�j�ܕ#)�@�]�п����R7�ٻ' r}�w�����#��%~:�$u�vi�0�N)!�
~���F�Gx΅�x�(߉��ՠi�ஂ�={d�r���"p>#�H-��1:��􇉏����M�4�ڑ!�:���zӘ�̥dd�a�SI?�H�O��g�-�M������3a�YNS�k(����ڶv�j�js�.~�������2#��xv�a�(s0� �4q�t;�v��^�I$��6�?���(1MM����D��~�w0R�{G�c��EG3�	��U�ev۽$�^W�1�� ���8˼�����q�J��L<ϱߚ�y�Ů}�pX��-p�q�t�]#��h�	�,й�?���&4�������Q!�{���_v3p1�<�v���ђy��ﰽ�ď��N�q��ޜ�BU<L��]d�0�ڑL�<��p�?H�2���g��b�(l�J	��ylq�2��:��`�6K��~	�5,Kb�I����Z3�)��F]b�ϻ+�;.;p�$9������:��.�r^�$�Φ=F{ӈIw �Yp�B���-��h�P	ޥ�hK��3S�����T�+ˎ��x�L�Ȣ�f��vv|X7R�-O4P$0�`��%*p�DKܧ�:��|?ƅ%'d�-.9�\�
x�'Y3�>�o�ㄱ�>k����}�钂�Hkj⫐��
�l�Dn(�~�;��=̓U��d���ZT�ΟNU�(@�0�n���1+<o@ﾊ:)�F)�J�;�TY:�q�<S�����L� ��ʲcF��i_ ��X6#�5AXU񅢗�ٝpಫ�q_���*��\MRB�׊HS�/�-�-#���|B�RB01���P�Y��[z|������La�ytJ8�t�b;��v�g/3�m�ތ���݈����h�&	?�FY��K���*z�`�`�q�N~Tq���Y$씟�ʬdGg��~ۅ;���m�I��f�4�s
eԮo�X~��y����gj��p����]�u~)3�ș6" ��*e��CK�,Pc�C���L�fwE�7���B&�
�N�;�Hn涂���BL�.gwS͛��~-���ZH���J�%��m���*��� ;�L�Ћ(&���u֣����JQ嚘��bQIk�Ve����XM�	6���|�*X؍#+��RB\06g	�ד���N�+�䱽��{��z���("���+��/=��i��M��r�6S,mknu��kэ�p�%��z1[��>��ko�~iv�DV�2d��㩇5k _�����,�eWe�d��!�S�}(�!!)�y���n�7:ҶZ3኏DT�	�c�*'�^��<���KE�r�ϓ���t�R$�(^�c��T�\n6�K|���o�-�t�K~���D�K��,���.���w���H��!!"X�s���).v	p��rH�]�M�?JD�M����I5�R�/����_����]�V�x��M&�/�&�R���Ny�@��g#r6� P�spM��b��������EyyDm�c+���Z��ܡ\�=�Ú�5�������T�>���N�G"��
u��� n�	R����)[��h3i3�j������=�7ZV�Q�	��;����Y9�{�G��J�{Ώ�Q�=[�H�˚�$7#p���ϻR��r� �����3W21���.7j�'�mA��b�����C��t�b�x�nn���dw[�@�MQ�,E�\)E_�;tJL���p��DY^�K��ϐ{�r� ,�1��=T32���r)e�	&����k�	&'����8R�s<�����j�^�= :N�j�$.أZ!m��N%�@�!W�;B�u���$/E�t�� &��9�ı.^��T6	1T�
���������-j)}�%�wp��BuD\N��)п��;�[̠��&�A�����s�
]{~���)�����?�l&�:C�\�3���y�7h��˿�/�|H�%����������!4�Бšt�t�f��U�%Z�.�|�͌� ��x��R��D%��"�I���T�M�^��񆋰C��ڑh�G���<$|���K��I�&�4���ۘ*,y���z�ё�{9��Ҵw�:�������+�[���Ҫ�P��F�`���	t}~��x�`ˏ=7G�2}͝��b�ώ��g���YKwR��
|�ٲ��D�dE���7r���D:}�7"��v~����N��L��c7�R�(��l�>�x���5`��(9�B� ����R��b�!yN��~r�[ ��:����mq �+�����g!�"hr������ha�%)�݀ޚ{�"��NuY��G�Sk��1]��ħ��R����Q�ɰ1I9j���	J�ۋ�br�"�)"���������K�[g?6�jJ�XT�5z�m�jڷBg��骷������x�Ʃ���h$�Z�m��|EZ���ԙ�*���9�l�>j�����ٓ�<	�h���i�RF���M�p�>+k/������l�d��Ip}�V�ه��3�.��J���IF<��W���r��rZ��X�|�5u���*���Zyf*u_@|C#W�ib�Æ�T����B�����+�0#�V���n���<^�����������Bp�L�/�3|`�d���	���5�h��[1m��U	s�	=�Qt��<��@<���`���֋��u`�5v����Q�	������&�S|i�K�c��,k�ؾD�E�U���P.�51<��`���_�V�AW/`�V���uch��h��:SR�BC��Be``��k-d���$>\������͕׊lw��$F+���Av�k�:��k.wF68�,�������'/���q����ksq��!\mO	���d�~�@�Bth�$S������E'u��Dj��a�㉖"H$��i�%V���XPj8���>��+����^�RgN��}�n:$��A�àݒT�9��O����G�.e�tn�p�����Z�@��q-D��~fI����d%,~.:�D��zP��׆K2�,����:-�6$�YAxP��h_��G��Q43���+���K��6G(���ڗ!����v-�i��}B�]�N=J���L�Ƃ�	#؞I�˖p��"Y��k�hsU�~�\�����ήg�3��H��T'U��c�?s�>쎗a���j��t��V���%lY��S���[�Oe�`�b�ٌ��i�������ÖD������o�j��[��+�/��4��)};/��	cV�s &r����~1���D�|�_�S�/�?����dRA*�AO ��!-dP�'@�Fcbӈ�Vo�̈́�6˗�c���JZS�:�T�=�uf�7�,�-a�Ӵ�S�4�.� �\�H���G-���-�7����ޛ���*��/^NÝf��	V^F��^���B]�=���9��t� ��=*��e� ��sQ�7g��kL���&��|�*q�︼���n��v�����UK���0�� �BƱ�q`��Rc�4(������/�dZ,��6g�7X���R�@����������áU΃��)�"�R]�I�8b�22�16Ɩz,��j��G8[��{��&�6N��bk]z��g����t忯@E=��1.ľv�u���W��D\�ޗ�]t�V.SLaLY�_��G��l��<Ϡ}��k�i��g� �B}$��u�7/���tVݶ�l6�>	U`���fuVfav4�w�^p&�M��z"��,Ds�k����a�3���6ȷF,�	KТ��U��6�(%�-PT�i7ڝ�I[-!����}�\���5+��g삷�_Ƴ"�;�MO{Ǝ
b���$�R�?AT���gK~�4Y�3'��-8�`dl�6����8|>��G �YV��k�e���;�� ��J�a'2*�,��aS��!����v������;B�df^��[�y@2'g�3×�9i ���r+w[��'�=\]b�u#y�DV^�W�՗�-�v�,xo �N݅��m�t(�`Q��=gp�D�=�P��+5C�&d��!��+��?�R!��v9nx�]�F���tɳ���{BTmm�{���`1�gN7 M'�`����N#���	�u�?��
�[�H3��W�����-�ܬG�M�3�}�4��m�GK�f[��R"��������ﭕ���x3}qi��>�+@!\�E�����o� >�4�8�{2�(����Y�h&��������z�筜W��a����_q^� yX�d[g����V$�7���зH�Y�R7Zp��*����5mJ50�F�e�M�?�Y���R�^�-��5K(��յrQ�G��KTb�;��g��7R�EK��Nh�5���d�}�p$.Xbr�0��n7�h�3�,5�X��@-;F�X�	�"Ӱ�;/���R=ʾ2��y�̕��2;���e�l���`*$� �6�Y]�m���BH���ta>�� p����Ƨ6�!ta��`��_aq]_�]	�+X��q�b���9M
z�*�"w�~�Vu�G봪܁���u~2��
���Q�����Μ�D�_��#���L�w�5
��	S���^)���Zc�i%gE��/�l�I���3{<��i�z$�	G��ܔ�-oc0�`� 3�p����8u0G��5�Y����3r�U��<�U[<�V������Įc����0�t�,��^��6v�)H�'�Z��|q�F�	Q�Va�l�
1MȽ����vAS3��B�g���g����(�����Q���G�Z]���;^pɷ�Y6�hw|N�z:�Jg�v��
P�{&�nsC�I&��z���;I7�!o�>�'�����u[a"h#)��2y�nAQi��]뤾�:{��K�m$��K���N�O�M3_�>�c弗5$���^H	�"�rWQ��2rᳩMj`���pCɆ������zY�/Ϋ��aE8k���1i|�tk��ˆF��h�DaC�����2���݆mC��F�"Hh�G��"�}��ߡ[��^�N�b��||��f��y��7����"�Ү�_F����?{k`ޮ.���1�Q=Ő$�ݹ�ksZ��hx;W�
e�r�-��N����`�33R�3�C�fPrPuk,)�8�l��M�-��᜴�{CVPq��Nw��	�ý��+ߥ��'��Xp9�kT� @��9��\Z��$|D��j}��xavk�c2x(��O���a�;�[s^�Տ��8���V|EGl�\eD����d{4���JI�p�|j���m�u2q��!X'�>atoB���\bk`.Q[�<	�;X�h��ٯ�	1�
�s�dؘ�~M-
:�S�F�:�{����ڰa���ǩ���� ����%�<�)q?�/��ġ�}�3�R�-��n?Y�[=;"%����!�z�W��<G�IEJݭe��#34\�Ɩ�D��m%{�ā+y/6r��%�/�OX@���6��V&�O6���b�#��:��h3�bn=|��*�#C�F;#�xl3�Z��^Ó���{ù�V̒����Otv1,�	�5V��b�2b��Rd�i-W<b�C�JC(r���X���0J�U��]��*���F�`%��>x�;�C��"q��)�&v�:�����z�1��ӂF=x��W�:�j�P�y�	}���Cl�{*^E�S���m^'�T���ԜAz;$����Ф6|L,>���oe8�,��[���68g���ƹ��b�;�jB^�����j1�6��;'��>�o�VP��!7�2OZ���\�'�܃wn^(p%g~R��yկI@#��qF2N:L�?9cM�*�!?�|P7ږ��Ż��s�F$��1�����xUĆU��ć���z�{���6Dl�F^��=�O�rG�9l#�31���0��`������}X_w�s�:6$��#��	���^ E8�d��1ly��(�Y-ÖS����K������~W~w�<O���%�L't<�m�o?��kL�Z�!#=9�G�z��+q4EǪO�����l7����ؘy�.��L�P.C�ΫcM���0����Hh=���T`7�@�P!�r�*�R8�:f�+p�J?��+4��m�U(B����f���̝ĉDgi��w6�}F6g]����H'��C�s����[ǝ:�-��7qN�([����L{WR����fV^��U�ZhE4�Mg,n�i��wY�L���6k�֒1��$��+T��B2�{l����[#Bzl�BW�z�J���Q�e�,�F<� \p�:�K� EڝH�v��f�_줾kD�K� !����=��J�o���*�}�0�]��X=r���u����	���������܃�F�6v�X���׮��u�4�rv��W�;��`8����1ױ�T�ZD���&�᠈Y>��M�����@q�a����4��։�M|���D<56�AcQ�7�WЅ?�M��t�Y�P}�~�9{���&c�,?f!�\�cc���U}�]�d����9�J��Rpז���=�?H�gPHK��e�C���Y��q����0-9�c�!9�tw�\���u:_��|��� b�gTɊ��'�T�a-�J��G<��Wv=������t�_w����ѣ^��Sl[>��Lh���Ր����J��%׋�B�{u�i����f�
��]���\)W>xG'�����D+�����yn]S`�E�\�-z,i��dȪ�=��ϱ���,bJI�!S7��`����[�e�Z?<s�Yy�+�RI�@�6F���oV�'�/�,�R�7�
�?B�͋2Ї�n����h�,��u�n�;D�?FN�:���F)�:���_VF}��膯I[*�w­��:�~X�昻��e;I/�&��O\xF��$_����>���vu��
\&�7���m	#p��_Lh�4�����y�}������I������/�ɣ���gS�nʉv5/0̑�>Q�pG�� w�O�L8; ���?
���f��M���� �?��f���T&zn�ja �n�T��zh�7л�rV)�yӀ��%/���j�>�W��:�ϧ�ZA��s�;C���uy�ӬX�n4w�����x��P1���/�d��	�:�0J�c(��Z���U�$ҁ��1r5������5\�T��̷
7�� �ħ/=]��4�-0�Ռx�֓M�5��D�)�(̡��X���.~��c~˥O�C�}Ɠ8:���m���C���*��TW��=�bN�O�A�[��i��۳��VEz��~*`�7�g^]R��Rߗ�N�2|v�m�1� Pz�0x�/> �f�2x=ޱ�)��tl��C���+T���1�����?���RH�S��+5d|�H�ޏh9[5�쮥ŢP�f�oՎ*%�x�;:�{���Gq�����E�3��Y���H������(Yn�	*݁�+{��-�uqZ{C�E5�������CG(j�C��Ӷ�!�fţϱu�[�	$�
n\!�E���;����$�G����5��r�֟l�7���0�໳��̥Y���v��W���`��Z�6�E�aQ�n_�G)V�	/O �H�o���Q���i��(�;P�柪��j� ���݄r-d��Է-nPvm�ײ��Q��J�����1��+8�H���3-{E�U?�g\_�\�
6�A�HDL�oVʡ-����UX5��V|���
B��ˡ}낺�u����0o��y���\���!���}Vt�I������ �}}V8�����/£Y��'e���~��:Kd+S�HTv�ݟGc�k����K�B'��Q���wIZG��Y�G�dr .#�꿦�`�:_q@�z�Z�{Nj&��������2��Sb 0h{�]Y�$�۵O����ٻk�P7eInx7���tm�i�=L���]tSH��':#�	���~��ubXP���8����
��h���|�שu���ufQFl@)�\�l�`�pv]b��`B*N4��Mx$����Hv�Z)�����m�*7t��^���zT�,{�k��|��10|>��-?��kJ�z[�ڀ�G�x�-	�2#M����dؙ�����X��@��=�ź��Nػ�!�N�޸�С�B�Ə��:Q���ŋ]���7�V��mѨ��V��"��s�+� :�D.�� z�K4��4~�O%9<.���XHn�y4�v⢳`�Q�v���|��$�E����ث��&vS���0BL��MZl!�7���y?��޵-B���FQ"�s}��~�:bL�_��jek��-�ǟ������k������Ǵ���"��{�(�_l��a����k:��2�7�����g�}|��
�~<�(\xʕ˛NJk�$��eD���o����Mg��z����*J�n�Y�x�g��Ź��LTBY6�~��1�m5���n��m� ��ua���%�5��a��m~�i��m�B|��W�5|���?
�����t�I��oZ���/�b�V<�J���0ޒ��[&�(yQ���Ao�K3�K����2a�R��%Bu�k�I����N�3�F<�X��p�]Nᢥf�Mn��B��b��D _�=@"zW��Z
aG����!��bH���l���4a�Цx� �`8�����"�!v�U��n1���w����l(���'J+�^nN�<���b5��7 @�����ה��7G�M�I��q�4��ŋ�!�8q��1
���H��P�_�֑�W����n��Pc���ZA��E�ݴl��1�qƅm����c�\L����oZ���r�����VjI�Jo�����;��P������xPs(�h
x�s�zD�*�}�G��̈�TLw�,q�����;�r7o��ӳm6ͱz/�t�^��R6�2ez�*/Ҵ�1�=e�\�7[��ɺ.��6�19�q&�Ӥ�AoY�H�;l�xK�(A��#�gy,��%z���J&��T�$�Z3Ե�][s$��1>�)��f���7�0��HK3���"\NY���Tg� {�"&g�2�-6�V����@� �64��u	�^��c�N`����n�B:(2��,6x�~k��� �>��.^��;��M	#8�6h������	y]����kO�z��Gk89�w��bu5�j��wz6�.�*7�E���>`p[���_m���@���/!�	F~��p�(�+?�S����� :�>��&�������11C���HGE^ۘY��Z;���]|�N�^|�yz�6O_"�����^�F.�5uj]%��ǹ��j�%0>�DT6�e��S%���G���<u�R\� ���<Y,G��."����r�����"èe�t��hh�l1�M����n���{,{�q���2y~ф/o�*J=/Q��}���,���)��<W��J��~�{�̸�N�8��$���5�$)��c�સ��Y6��fB�P�u��%��f}eH��E-@�����ָ�B[�� c���n�5���/���Ly8���l���r���_6��D�O�%��������G�0��X��WR��6~�����������&�7Y0���gE�K�ڴ���Ҁ��r��cT�r����##� /�#�S#���\�����'ckmjK_��:���i\�)|��(�^EDs�s��o}NZ����nQ��w�Anڵ���������%S���H��uq�W ���G�T�!����L�7lƦ�1!k���i�ń�9uT'lY��l��DgN���W������F��P�[��n�%A�!�W�����j~�N��	=�#3�%�k �)D���]�ƒQ�+)c�������-���\OYi��T>���nݼ���7��3@ (V-3e�.� �V6>8�v��G2�f�尡�c��,�ήa�7�������&T�9)1�c�h��񝝁�Ǣ�УT�%_꘎ �o���Z����������NN�\ҧ��F����L����ӿq���d>TۺF��mG۴��������;��$H�d����q�Z8��5e��4O���s�8���kWDS�넅�k����G����O�k�AO�K5�f�Eo�>�Y��r52z�6ӎK0i��.(����R�Z����s�z�f����{�N�>j�������Y�,dW�]���q�II�r;�U�Y��ŮMP"h01@&�ْ�s^5R��,�c/9&kUdI�s��-��J��%5H�/�#qI��56�Y4�>�74�ugMq�1� �f�L+�U�,�hu@����`��Pi�)�ɟ[]�\�����f�����x$�3`��#3th���+~]������\1�z��"pGvI�
--(>��
����\�����)����Q��m��P"^Bu��1��|Jt� B� �t6��07����n��]���{m���f�(J��9������C��J��y��e܁W�v:ݼkZh�S��z؎��v�y��=F�\j������/AE%�����X�:!XQ���TU��YV��� ��ra�0�̜�MP(�׉��7$�ݩ]�v�LPf�z��sE���U6��p�b�֬ݾb�+2s�9K��"��K�Q]%�������Z��;�+T�Z;��B�P�n�ZUb��{�Τ1K�|�鋅��	�"���Y�[����D����N������U�����C(��7�
�-kV����_���͕"MF!
�Yo���V���֙&:u��h��l�RA)�F4r��Z$��8G^��KTr�2bĺ�$�_<��'�'�|�����h8&�bQg�V>�S�����1
l��ߤ�͵ð#�M�}��AX �@6��[5ۅР��_��8��j�
��?�W�L�u�`�8��#����(-�9�P��j��c��\kZ�~2U�ҡ�	)������Z#�:�B\�-|׮T�T�j���=B@\�^��s���X�����}ϟ��$�p�.��L�k2�*� ��}���u�OL�u��j��s�� ��x8��ze:�G���n����������!� ���!W����Ok�O�
�8¯�s��Dn������7(������F��������5�Y�l�w(�>��4� uxm�E��Eԑ�|M;3{>/9�р���P��g V�顴�"S�L���|��p�J�+Y�`So�&��n�@�"i?13��U�������)̤u��I�p��u�o��;��*�j����N_N�d�
�����ENr�;Q���0�$��con��0�<l�	E\��;-@��.����S�Ug�T�;�F8�L*~5-���[{�@���߮2��I��W-�inIK3V_4��>G�cA0B.R ���X�Q������)�4�{`�<ty�����_�A�k��)�mlEDG0��?��bO���WͅMfO6�7��Jm�Q��U�t��׽�<�z�	a�[{�����4��k @!��$w�C?�u(.뗶6%���\ v��f��u��W�
�4���{7��h� �*��'6ţGn�����x�m=��[`U����Xb�9N��U �KM1��Z�X�½u�s�&��9���0�Ƌ���'�G�zK,���G����GS{�v��/wg5K���W�fK�C�d�{��޷���Z�&�L՟���u������]���"��\�c�Ү`�(v�����Z�mtI��4j�rѠ|E~�@Fƃ�tT�C�T�Kȏss+9s~j|1�Q^﮵��q/eB.�B�!��?�����i$%9F���3>�=��t�U�Z�q�z���sd��+bڙ�"`kw_��xF�o����aXuD������q���B�0�l��It:Tӧ�b�ȧ�����y���HsM��R,�j�M�-�ߧ��ZZ���En������� ��NE֚ʺ������ ��h�F�]ݕ�ԁ�{�ԇ����eT��gx�D/��o�'�D�1&^��.�|��u)�rc�_SW!���*��ra���̉���"�JF�@<����O"Bl�h����q���Wy~jgjJ�0�A"6�;O[�Y�����Gүjq���Y�=!�����6+nNR�,�N�l�����;�����N�J�?7�~#V���թ�f���\��}B�W�O��?!h3!�U(�l��Z��`B$�1=aҘA�F[�\��.}v� ���-�c��T��'�^VpX�L��K�>B937٘�~��QK��&�`�!Ď0�4���w�!>� P�B�7�c�qZ׷e���0����\xC�D%��JA�gl�ֲ�-�a��'����I���h9t�#U�#�:���k u�Г>4�q���~rп:�	Ȯ��u�(�T�V�<���&Qi�Z�B��^�۰·̘;�_b�:Fk��Tl1G�!�q	hu��$z�����F�����-�W�̽p��s�y�?U����-�wTD���ve,�U
��"J�А8q�>mp��Q�XzRB��hK������C��� m�r�_m)�}7��s
�����a(BsJ�KYz���S#�/A�5_��q��R�=?�D������!�Y�c T]��r5[�ƎJ&�[�b��)g���0df1���Vpo���x�{X�L�j���
f[q�N�v��*
پ�n��⧒�"���p"ߣ�2���u�}S��`f�eЄ� ��D������8���9	a)�i8K��	R���D�������'��X�Ix������Ԓr�Nt1��ډ|��&����G�� �67�+-@�����3&-�W�8F`���R?���������DQ��s^v:��)��7��5.	�̈J�2��q��~3AYU������-W�$�Bc[��P�m�-r�l}��7�v(��a�T��&$��DYen<����>�E�� [Ш0r������T���0��+������.\sa)\���&���f�.�$�ӡ���g�U��� &W�f%�ɭ71����(����a|��Me_�)�%��j��'��~ݲ�n����ǉ��0�Z�E!8����_r���%�<�{����� �U	��L��c����r�ΐ�hNS唹��T�8�8�d�P!�ҭB-�V�ª���<�@H��^�#Ǔ!�Sw��yY��P�C�:���>ނ�?&��w@e��k��{J7�{�V�G���e�	§=2D����5����֚7.Xܰ�Z�O����)K����z�{%�U/p}L�EJpX��	�b+���������:����Jw�Y�V�(�i0��Ȁ�c~�u	V�s��9#A�y�v��g%dMe�:����Q���Kxt�,+�Vl���lT������,�Z	�qW��a��ȝ�Uh�.U��D%�-�HF���܋����H��X�7��J�c�m~����X��$��ju&%=5F�?�Ӝ����+�@p�$)	*
|�T_��Wɜ�1��4�8�S2���<��#�W�<6��eBGvsß=��f@�nQ1��r�\w�$�LDgO��҇�*�2"Z��hl�7
��W�ss�DDe];�t�9�t��Lʑ�U�Z��йS'mR���s�'�$^PmR��kB�wu�}�eP�	=�^�'�2�-pu"2��JS�٪OT84��g@C4�����s �4D��K�.�o~�H ;���;ao�`�����n��{t���m�Ѵ6x1��'��\L���� �ԁCxS�me�)|t������{�w�p�T5 ���NK/����-��;|�7�*��������~�M��W�ar�ԯJr��nwVF5Ò݂�)A��R�6_���d�N�A�T����eanM��>M$^�[~�XG'�?.6С	jc2�]��3�Q���H1���(�L�.�`p�U����P��nn�JA�uۑ��וڂR?��5��\ݩt�c�B���YX�0�0y���X�5�i Pc�:��k�㮱W�b|�-��Ԉ�ֻbm���6���R���j;�����y##���ߡ� ������/a�}���jg�88������¼zT� �5��nq��i�Feh�՗(���~U�0�/@�x`����I���<a���cy�M�3��f�����)��*XQ�K���r�<*]nS�3���`V&�W���dbA�Ys��X-��5� ɩ��v�l��iV&�v�0i�	=����.�
�M�1�M��ڋPz�A�ۢF���ⴟE���7���(>e9;5�g�$� ^�3��c��z��kJKnXr�r�3֣^������e�\�_ꪤ+{mM�������mj8�VnE���-���<�.�%g�'��9\�袋��nX���C�����kS܎0��:lǺ�v��L���i�j�.�4&p�.#�Ǩû�3��Z�[{�eaZS�-��o��:[��$>�k#��6�v��GD����������݈� N�1��n /�����DAq)6٪�v�чӊ�f�qh� '�2*D(����"��Ct��a7�{@�ͤ�C�hvA���Ū6��t(,ԥ$�Vک�fуY�TpYG��T&~�v(���%Q���|���/q����%lw�m`pb��.���])%h�. ����UPE<�i���s� W2<�*e*�ô	��ܥ���U��$-ѫ���@��{㧠w?����j�F
?�/�Dqs�s0ɶz��3mx%i����7�CSiB��XC�τ�Z���5���tH?g�w������	i��u*�a��W�����̭�L��Hb��K�I�hq]�����(�q���AT�~����m�(�W���?�������\�oH<�Q�Qk~<+�=5�-d�l��v|���݉h*v��\-"�nR1Lv9hg3��/�=��)���~���%�[O%x���Ċ��'��*�J(q����� l�lu[�����4��e�x���3<!�k��T,���͡bkpLd������O}I��'dw�[���}��E��˫|�q@�䌑t�tU-Go�c�����$�K5}`���H2��OO _����c�8�ɇ74R�/�E{�U��
��40E;��0G~o���l�Z�G��k�_mCȽ�A*�S���z"9����Us����)+����G�I��t*.��^t�-f ��rbd���gҎ>V��U3�];<v\W��>r���W�OŐQW9F����n�+�'|u��%$���}D��J�D[��À|t?� �QtM�;��ߔ�6�rj�ٖ_�c�	K�i�o�Z��*�G�z3T��1����MB���A�	�V�	-Ȩ}	��?��iM�@@��U�ץAW�,ק��qO��Q�*�Uǅ��ɍ*�����N�b��~��.�m�3f�7���4�̫kf��Em��Y�3`練�h4\>�G(��4�&��zn�ڴa�����4�/3�hV�E_g�o��0~��i �&�'�:��j��^L���Ge���E�p@vt�x�Z
9A�d���� ��U��l�Pz]\���d�Ã�k��m3ӱ�I��bЈp���e�7�MC�}C倚�^���we�P�~=���.g�Z�)Y�&]�x�c�7��r	��f;i9�Qn����܃�^^��ڢ�L�}!|��|8����g�y�F����К�bs��Z��<�S�P�$�cVw`UO�Cj�� ��i�"A ڈ`d��q{:�󹀒);y��+DA��paE��CGɻ?��_;d��.]�B�L]A�[������ i����L�J��'��IH�J��O��@>��ScV!_i��;�l�ۛ,zyw�&��bj@���T�cG��&���:."H���+#
\�\�'�r���e�s<��q͔��.�����I3�돘�}ɋ�q�-�/"�����Uo�9v�ڦg�*��*�[��%�_��H}�0 ��<B�*8�c�W�g��,;�Tpm��ɗ��GM�u��&��y�rB{�q$�?�_��!.�"�j�<��g[��&j��HR�u�6���EY�٧��+�9�)�f���_�s+塱���@�ҵ�G���8���1S��90KJ,D({�v%��N|	�&/����q)�E���c��p��S�i���0WP��"7]\T[�1�e��9���}YPP���.�ًk��{Q��9����@����ɰ����0�'�*�)�S�J�͟�F4��1}"}�:�]Q�r�n�7�m]�z�ڂ�(>:=��ĩ0�XoEzt�.cTˎ7I*g4�
GuovY��Kir\�i���6i@��2A�Pitʍ�غ����N������A��QN��]$̹/��54tl�J21�GD���wT����N�#4����1��7d�������4�lv���O�{R�| �R� ��%m��)�*�+s��N4˩D�6�D��Fz��L����ź(i��QJg�t�4����c>gmexI[i؁\r��"�N@�OsQ���qF�n��R��䃓�eߩ�Y]yAtr�J�_~����z�_ڳ¸s��{SC�E�h�,S�����U%��X_��/���~D;j��k7Ü찎�{�&#o_����L�{hpm�V
�K�V@h�7Ţ�wO�ؓO!��\���n|�9ևb@wC]�>z�>׳ z��ߺ*s�X�޳�sk\�]�����w���h�c`!�I谺Orϖ��=(�;��s�V�_+M�@��E%:�|􊑶��"0	�����"�Db���R:ə���u3i��p~]^���lRPs+��TD�!>��T��CMJ�7�'KԟY���������r%D�Oa�3�֖qRh�N�[�P����٨mg���@�[ �z�	re������C�6��N$����DXX�eV���\�����A�UJ�噶����O�q��d?̿�MY���M�H���
\�	,oP�=G��UXpb�iQ�����b�z%iۡ��u�'�to��ʘ�2�d}����_���D��k�$�����i��b�X���)���pֈ�K��ԧ�y�X�y<�����!j�R��vX^����o�A�lI�f���	Uh1�_b�I�)�x�1���\d�zi����	o�X�q`�.��T�6/�fu(_�r�����O�W�;"@&�Εr1�s�,`'��Vl�Oǋ
�����-!|D7���@��i�#����b��x��\���B�N���#P����#3����~�.�K��e��=���A��EzM �f��g�����������Z(��ƪ6��*�N-eXM|%_��[!��AkCd��A�uA��xfC�;�iJW��G9 �A��	�o-��>Hn��s���W�ֽ����u��I��8����@���Rm�u(ₘ��*˄Z�C�J;�˼P��hLE[!h��}��'�g�z�h��*#���w�4Ӟm�v�vs�fC�3'����M�2��T��?��9B@A����ٻ�Q����R:/�@A�M�?M�.T"�B���Xv��Cc8zϕ=̋��}z���Ve6�ł3a�.�Ͽ�ɱg'��Rf�&ʂg�@�� ��J�B�r {n'`{.o[��Ʉ�(�%�`15xʡ,�<���x�]���AM�����N;7�}��S��b�����ҵ�X�L��S{�M,����i�c� �} P��I�^4J.()�]�\�L�	�n3�@����]cm�C�Jm(�S�w#4$}�B쭐�w���K�	1�[��	��wc}_KL�!�o0�%j�W�M��%�A�.�2$d�$�HoaI��0t"��&�!&��\����<��}-G!��L��Ԅn�f7�bSK�x��ؕ���눰��\�2s���P���L8�m�Ý
SxK:$5�N��'�TY��ϫ2
�ɹ�d��Y0+��1s+޿�
�
�/�CW7��@��@;���.��^!�6�y�������`.-�#u�Z�t�Ƭ������R�X�%օ;���T6 ��?t6�ߵ��\��y �4���A\���qsq8�o��k����籅o���/�)3"�Q�`�R�2�����\��ҵ�ʙ���4�>��˂���J��Q�Z��٢i���'��e���ʫ�N T���w��޽��-�2��r7�B*�'��|��/�jyLMζ���E8�j��!I��̘��d[�����K��Q�
�Ey���d�Q,�n|̤G��n��zP��俸��l��qqt�cf"���t9O�Z�c�ylJ>lMwMRpWۦ�%Zi�rF[�\��iW��=)���<��㨪4��&�בS/nxlIKm-V,ꁮ��STd,�U�T4C��L��z��-��7�H<En��m�oDL�Vg~��k�������f�ifߏ�X���s���!@V�����G��.�q�M�+�T�E�t]���T�ެ��*�i���PO�����D�V�[�%��\e���+x�2�%��d��"A�Ϫ�^��ł��W[� ����7��&C���:����&�w��rV��"��G�B3���X͸���<�/�+۞�v� �Ђ�?��}�u�ò� ��1;''��<:g�k x�o{�a_1�c��2�jnI��[�\��)z>�)G�,.h�`�� *��K�����{td	�Kiu��hZǡ.�V�D�����'L�*e�����~wj=U荫rP�ڪ�f��-�#kCf{_��ߨ�
���s�| 5�IuȀ��^��Z��8�|L���\7�=���O�+YF�'Xv%��pS�F�]�©>�ؘi99�}7 5%�3��^ݭmc\T��$�`� �=*B%��Ʈ���r�9��X����58	�"�~b�\TLv�(mha�Z���0�K���.-�S���^�U�7짭���D�E칤��8E^Wα���O4.����6��z��s��ׁG\�d]�q�|Y���ݍ����F1K�9���=�}��Gb���;(��Xy����MN�<���ܲj@�*Uw�{�,�Y�Т\�>�٭k"ѧ���$^��C�֡�̙`�Fka��!J��@�@����@����PBuO�6��8�}Q�0+T�1���ܿE�(G��~�{�C�э�e8S�Ƀv�8�6:�,5 ���Le�73&(T u�s�;�u{��{+X_�ֻ�tz��aa��G�'V;@��
ʪ�7������������CǐY�y�n��=���c��嘍Q�깣�f31��<*G�\���fT"ܴ�;�����A0A-��=+�	��^�E$Z�u���F6Mp�%�R-�gs:�P� $zGE��w[�����.�˒��xC;�Ė�&��=�e5���j��PtD���FbåQ����˅�V�Zܘv5�1�f�Y
�`�+8^mݯB��l������i�c�x�fE2BMe����r���}
$U��?����;��=f��;N�m�u�����*�'�<������ ����(#���Lc��AvbpH��!Qo��_}V2��C�~,Z��g �m@��o���tXY�Q"s��v���a���-�0})��X@G@�{�^�vک	u*�w�	N��g�ƺ��pA����z;W�*y��Ln�J*X�����P�Y~�#���ь#�޿u��e�m�_��ޟFp�U�T�M�0�Y��k?r���n����ed�m��{��;%�}-c�1m�-'f���EY�{:�@%�mk.BB�!t0�h�2=5��I�4�z��pVo�ҝ,F���,Z��$�'�@>�G�"?��ɥum��1��:]<�P���V�W�;�lr��T�|�E��!�W���W�,|��-I�_��^3l^�.�ҍ��2A �!�{���a��ŵl��x���d�9�V�椟���{�DaD�ߘ � �������~7�����:0x�4�Z{�Gp� \�J�oJx7��+��sn�
�% �UnPPՓP�2�-�7�QD�ԙ��'Eh���$uD������9D�Nf���GVm>�����j}�n��zC�M��4�^X�@a�!'^ʿ%&�k�F���-�Y�Y�T����s�c\�;6�bqYe]��h�3���L��R�y�O^
>�����-�S��ޭ�������h*\_h�%]zl�n{�6�Si��S��o;������ŝ�@@�k��V�3$�\�}w�)�Hq���/�M������ED횟!�	5�n�j<�_���'�M�C����s��W�G�+A����}NS�U�h����P8����𔛮}��?���쵳s!l�*M�U��?�hp�"�T��h8�{�y�*+Y��k�����XK�����`u�}�{҉��3��[�;`-��0��}��*kGkG�U�$�cA�
�H%�y��u(�g���`�$�8-�{������r𹑨��-�+&W{�Ѵ�^K���2�-u{��λF�d�4���Q_7��/�"(�N8X��>v�u�T������ �J���H����[�]�bHg�A�E�'��ԧ��K|�n)�A��,�c���v��hT4�2V�,�������A�f:e��\���|�{�K�G�l�g��کmc�B�'NeB�}�QDB-=�+�䁔�|mݢ��pl>i9­�'iL���mbt~�1Z rJ���0������N�6���K��Ȍo*��f���U��VR�D�y\��A+�_�-e�d��B�Gk^[��!ܼUZ_��ވ�Ź���}k��v���5�Vx��Ѕ��#'��C)\�T���7*�+��^��;(qLw)(��X	\��l��=�:��f��	�ю���p���yl]��+g�� `�&�Z_�ܵPA@�"��Xǚ��D�V�5�����
�ک:���ĶJ_m��#A.z�}�?^R*��m����%b�"��*���H_����y=����9�{���/��C���D��m�42�%�Ҍ:�uԧVXs���5���>�`q-����e��i� �ج�?A��@�˅���֧��v�q���a�'�Rҭ?w���ЭVm�$=0+�G[��j�p6�vF+�� �b-�V벜Z������4FǛ&}D�N��A��P����u����;`��[�Gv/��q�=���{�>YE�(2�?�=Ϙ@!G���^���Y���Z�aZ�6�V����TCu-H鼿(�g����E�[JcV��;�$���%H_�vj��{/�;Y���x ���M�"�r��V̵p9���_~�	8��L̐h����Rirŉ�ւZR�L���D��~*��B�tYX_��iŀ����T18
]�O��}����x��GS��b�|,~k;h��VP���<�*�����_�x�����Ik��3��H�"��R�ѯ��vq�����w�]I�2��G��X�13�>?q���w��_�WY�};rA���眺��	�����!��e�YoM�W=bL��~.Ҡ�+��k�v)FMڸ���0A_�\�6�������7�O�
���&]��ceYj(Bu�Lm�Ai-�LJ�����N5�3�	�0,�2ݒ�'IF̀��Mk`@g{9�M"���iҰI�m'�	Qݣ�ǅ�U�KB�]\�]�M�`�5;OS�w�����x��Pћ�R�Hp;~��~�k4��� �T��y�x�sL�z��?�Y���~Y���og��D�>D�(D=���zg]�!��N��ӟ���Ǝ�~'����3�*��}�G(��\�t��� ,))�,���wI���������'C�D~~�~H&�k��%'�ڜۈ��8"|��!_��S�l+�������6�4ï7��|ʮ���11�^�"�>y�E�L�	����s�� ���V��9��Õ�&G(��H�r5x���2�c�Cu�Җł��i�"��:B���}nS�ΰ�+T����>�h�n;@��pA�� W�$s�u��e�^A�%��� ����i3��!f�`4e80��6d�q��������B�S�9�l���=�^�E*���zeS�:c~%��8$�X�aV�>�0_���l�R��V��L�D��6g�E�k���5����+�L�nr�Y_��l���t޵�"�}"?]���F�#x�RI����X:U:�@�q�b$�J㤚E�6"Q�o��V �l�Í��	%ʡk�"�b?Jk�c���	�6��R�uӽ����5m�p;{�N�z��F��̆���RȻB�t��`cW����!91�~�͗`��BF�!fFC�����s��k !��J�L��:��kH��8�D"^A,dI+�qb/�� 1uDsG��i�w�-υ�w0��+�P*}����^�m�4�A���0�NMůU�`����'$���&��Ÿ/&D)��\�T����F�g�Va���j�"�I��P�F�@��
W�ׂ�/�B��"�ú�Q�g������>q1@����e_���a*���~K�D�0N2�/�7�ҔBV4��� ��R���-���/z��t#����4�?^����p+�����W�a�6��ܲ��K�Ί�c	�@{8'������/f�o��G,z2��^���nN���� Jî��Y���\�M2ҜӀ�q$$S�[�z*b��X�&w����E�{����z��*3�Cˇ��!���}�GY�l��Ÿ�Z{�r�6OP1v�!���h= yu�r���fB��u��>�Ih�?>^�1���ƶ�Q&of��
\�3-�]�i�mֳ�� b�*oQ��Uɲ$7b��W�{��|J��*�.[	fa��=69K�%�h��f[��:
�\�th���������x�NA��d�\
��L��
股��w7�ܦƐ"��'��îɽ�h�N�cղ �ף&��4�e��F���2���^�+H��װ�o��f<���j�3�xWՏ�]���� �.�2��C-t�Y(щv��c�4�:}����V��/ۅ�
G��	U'XI��N�o�V;l�'	��Oˑ�m��Ə`��s��M 1k��&ч�1�E�k�FT�A�v�N����=�8,m�6WI�g��8V"��Կ�%�\��C@᠅����s�A-V�����	<A~��Y@���O^�B�08)�@�a�t~�1�^+�#5o�MˮS /�c��b�����2���g"�I�&�w�$K,��<˺ [z�OL�T�')e�f�qN{Q#���/s�$h�T"����Y����e}7�P�.KG�� ���Ih�֋��
&F���W=>���ԹQ��s)��7�|�����4��[cd���d9�ٮ��B��M�Q�3�̔r���d���Seɭ��q���t�CgOV?��&u�!V#�>�$�x�*��ip��?�I�% ]��ײ�GF�Ţ'a�9W�m#&C�l,֛�7L���F��ŪR۝�K��&��ROnv)D���do6��.�����{�]$�&h��:�d��*9�̎e���DT��������<�-oT��>B��uY�������~Ǌ^��O�2�wl�-d�hǣ�m����)u���Q�G�G /]I�� )�0a�=И����L|��f^�N���<���f�;hԥ�?��<G���!2w�7�mpkS�I�d���I���~�by͒�g��-� �Pc&�i^?�I���J�J�Ƣ�r�5(b�S�C�����I�.�����J����a�!Oa7o�}���q�G_���+��m�� -�� � /���mP��'Ql�U'MʻMA��S��?;�8厕�a=��~8�#�V�ԩ&k��
�� �_�f#p]�đ�W���䭩w�^J�Q��	��Fxi��QH�{.��5��q�h �� ��{��	hv��q �>����S0	�Q�� <#�;�#��=�d�挊���x-}�Z��ReY���xE�b�9��#<U�O��'�l�MX\�r�c	n�ABݤ�O;U+�pq�@r�MH�c+a�Qdט���q��KwWk��y��#HS����E�=�
�u�"#�:$��$��p4�ʳ��RpŸ�+QZ�M[�������r�ˎ��rhRl֭wt^wshʕ�U��ƍ)�2�}��Q7�������
5N���.*h�bH�N0G�t�c�&l�_J͟��a�۵	=1�2��6MZ�3)D�̭b*H�?�,
~,��,�'ڙ�7���>|�;�"5V�n&�`+����s����+Hc�{�������U����b�t��a|�0��O26��a��oBo���3�j	�w}�y�g��X��M�P/'%Z��VA�>s-�(ɡ��@6Ks�1�45��r�Oj$�;�l�̎Zb���ꖎ0��Mʠ��|��0��UG~����8�I���݂��ƽ�J�)j!��]�^z����:;�k*�b� т)�$��U[�ogh;�c;�U�j&[��^�ԯ�V���r���WV��9��S(r*�����)xUFI��Q����A���*QG�����z 8��BYz��<�?_�1�r�V�_C���Z�AK0VN-W?�db�ƍ�a���G�%���8Ί �I9>n�;%�W�z?��!R�\ǈ�ݚ�OV^r�#�i� s��N��GSS�<oZB/Q;�(j�Z�&lUٝI�KkT�H�q5�a-՗p�� ]��t9��ybNF�:�z	��F�J������<v�&b���1�r3�ĵP�^���A�"��
c��Uօݩ_%�jyNV��Ffw�S�I�~3��R�f��믚�MQ�h(�y��%��G�֋�[Zx�bS�y�x8������S�BYF��Q��&X2zԈo�"�I�Y��k������ԃ���F]peX,���Qq�E0-�{���Y�W�T��w�,��RG,H$���1��S���\v�rz��=�`k��˷�D L�%�w�w��u��N�a6)M�"A9�,Sg,��dB=�̎�# ����?�0��y��IK
�2���R�B{��m��a���7�N#��0D�T~���^�*�rX�C�S���� �Q��Skj��sĭ'o�����j���|x���T���A���	��@�����H���5Y�!�zu����p��3�b�K��Cѳ�#�F�`a1��[�����g�W**�OJ��AC��1�>&p$Ϩ/�A�b�p.�I�{�����ܦ�����G�m��h�ۤ������(�9
���R���j{��X��;jr�ҳ���a}�Y����h� ���CI���aM��-u	\g*�#_S�w-1,=SR^��ŘS���g������\��^��KtWF0����c����#�n-���2Q�a��ײ6 ���ۗ�V�u�E!�cƤɍ�Aқ[/���8p)�eq��K`�	���C��*N��ΏbPPCC�� LC��bd?�]�S����(6�!2y�n08x���F8\�L^P�~�����b�h�����۫�y�_������u���ޘ=����da¬�A�}����OŅ��=\R��ao��(p67�PjֹLZ�Z�yl��Y�E+hꍙeh	��V�8������O6��z4��S����HnQ����)�%v�8ь�wY������MͬU��dV�kX����q�&�i��S\/a�f9���Du���#x#�Ŕ�0 �W���8�AW�8�@�`�8�")'�j��V����jd�
O��!�B��w���k�t� ٲ����^�j���s���o�J�
����]'�uV�#_T����C���D�Ζ�5k�����C�(�\�Rm�o�{8/C��� �v\�*��G��!Ŋ36����AxfOG2��m���E��U."���?w�T�Ӭ³���gߥ��Qhm����6�84��n��V�'��l�h7���k⭾�����	�H�j\g�㇉Y��"՛�������9�h��zQ�e�gl�]�v�藿ۋF[d�o:~�H�C�uTJ�8�W��{�~B���
��������Ɠ��ԑZh��m&�7�/��jk�=����w�'o������v����@����Q³-�o�}o��"lW��`}��5v/����8�wÀ(�N,� FdT�R���Q�"4b�/�fg�"m����FK���)��-�K�l�ll��5�����(1J�##���h��S��_R#����x�r��6DO͜�%8Œ}w���$�7��������I�Mg����|���X����*��(�%b�t���8�c�{����z��&}'�-�����O&��g<�L��g<�ஏ���G��&�ڔ>r*�.���Sn�:��&Vj�����Gl�S�U�,��Gb}�!�M�'C��(��P(�� ��`;a�#�j�����ɪ�JX�Ўf�(�*=��s��fձ6�RAm��p'G`�0��\����/Җ;�j� &�۟���=&V�jm�C~B�&����v�$�#wh��(�Ȋ+�ޏ�[�ē]����ԔWq�!W:]�e��j����z@�*{�k�U��̝dgV�4��[o4��5W������p�"(�Y:�a�Vo/��5��Q��٢��>*P�p��,���U!]��㋕��×^A��D(��+K�P�)�q�l����r�z_�m5��|Ǌ	/��(��[���<�F�!�tN����G��w8����?c�2�	;Z���{гSo��2 �ݔqCm��t넖_�׳^��d�o��_.�Q
�H͗:�l��K�?`���/V���kk,<}U�-�W�]�Ԍ4'*��!��;�t`У���}�9�s4Zf�+'V_��̎
�Jg�{��;���&�T�2���%x�F5�U҃0�Te��B�!�Ŭ�����,k+Щ� �:��l�	��U���s@�� ��@�y���bP�����?��jc7�a�OsA�WyA�G2Wz�5�,Hn �m�_z����Z0Xݏ(�.�Zx]#q5�lĎ�o�qd�g��[�}r��-Ow�M�ʷ�ٛ�,#��t#��1#0gJy�w��+�[�+�I��z�ª?��1�l�u��%jnLc땶�d��BL!�p�:ꂃ�r߆� �����m�����ꔢ"�J>��׫nҧ.Ҿ$ժ�! ֞��_�R�h�LiGA�yqG��~�x���c���ޖr�! Eޓ��^��t� ��`�g#ѡ#
8(��j�ќo󉐨F3a�@���$�%ksp��O�f������V�f�S�ҥ.(G9�EN=�{d&�2=x�R�v���iΞ��9Ѻ��������_g��@vǭ��ېY�hM� �.���h@^(����x$�e_`����EQ�2�x|B��Z�yQ�a�]/[;Q'
��ۧe�h����yp�����zL���,�8j�Ǭ�/L4�H�!��톐�Li6�_����Н�g��>{�(�j(2����n�A�'�Y��/��>��4z�bc龶�����fe�@�����v�m����h*��UO� s�=�ߜ#��14��՝IA{������o?��K4�a�;v���p�3V5-7�O�A��B~O�流�U=�$��{��{��~������J)��#��b%LU��Y� ��1h5�<�?�E@=��I�%��@�~��FO��^
�ƈkXq�B6����6�M�U�����vq��B�2)v��>h�X��x�������c��R���=��~�Hz|�߈`���"{�,P���5
P3�B�\����p_�B�u���E�(l\��^��u��]Ki���ҹ�M� T���;a�^�W!�1\��3�ƃ��ƧЧ�q��-���2Y�n�_���<P�Yr�i/kH���j�1i�h�ʤ"$;3m*9UCG�{��{��j�R�O-�%	-sM]��poNĎab�uէ�б
����p�#rY����Xu߭U#ri�|᫕+�w�WZ[BJ����KLM��U�c̽���TA^�J�v�Pp�;�=��� �����`��Nѭ���&����r�t6p�3S+��i�k�M��B>`U�͕�ޝ���~��\bgi�}�l��"���](\�����V1f���.��g��T)Dw���P����Ћ�6�P"��
}o�)�A��ص������pqF
���	��d$A���_nn�J�ڧ���i
;��O�x�U��V'�]�i�_��g;���𿉒=�)m�ʋ
��#����)hg.�bC<�9��AR�����X���
��g�v���/}L4���F����1z�`�H�uXfi����s�mR�N��e?������p��epb��z.)���OzgM�x��󤝎�N����d���j),�Sgu�4Ȝ��<�>��.��>1nh��ߖU_�ׂ�k��6[�W�����j4�2�����Bd̐�EÎ	��$��z@�)�9s�p��rn?�Di�/'<��!�j0��!AڲX]�6���,3��@E�c�7Zv"8c=���D�٪�+��W�Q��g
i<p.~P7rHw��6��7/~���2/��	)�4��R�)�}ƅ�RǴ�������(M�#*�/�_�rK�Q�vU;k;���v��cr��/o�^��Ⱦ`�u0�{�szkR�)���V$R$�bO���˶x`D�<ľ����Y�,i�I1|�t-�c�0���{oMFG	
�rQB=�0[_��ל��#�[�M�tp��!6�Dttc��Տ�>J+͑�*-2�ҞY@���9">���倕<^*��cO�P���7�!Q����L��>�ʷ�^�xq����������������+,yu���[l	T�h�$��S	� M�[2&��p )m��az���Cʑ��/zF��}a)��+$9��� O��d1���!P�9��_�s��hx>�H������a�V�i���,��Tl_�AeR͋�s��6��>���{�K��{���;�� ���Ο�BlZs���=�\u����A��s5u���0�@!k� �w�􆱺��^�x⊉Jh2��¹�y'��V\�=Z�|I����BO.�1��'��GaP�#2��R�_꣓!ت3Y�ꔚ�]�|̂{q�w�z�s犷y��J�mX��}��_�1��جB{��<0'zah�_~`H�X�ڰ����BS
��2����:�6y�*V��hu��7�CW�"uK��v^5��ؠ� �GE|y>{�+M�.	Br5F]��Y�{�ȝC���2����Iŵ�i4��a�.*��"v��*A�p~$M��CFk�p�fm�&�Ic�M\;ǒ�?�Uw�v�^G�h�9)�"�"��f)Wƙ��
��q���}L
�@��3�H@�e~�	}`Z��>�֦�	9V��m)B���\�5�֨�K6^h'{�3���ʿeX����h�W��WL�A�ce�G����� ��J�п�t�Ֆ�;�M#J��ZD�fF�*k:e�����)��B���f��q�ڜ�k�8"���>�x���/�}��<7��D"�wOd7K79�f_���g�HZ����f�U)ny���ѐ�?��&T�}p�0H��6ՎVz�P�2�2�*~�	�=8�9�x8���V���o�*T\Y��a�L x�|�F���PR�R��H��A�⁡z)a��s��I��ݹ]BMd�2a�TS<8��5-���:�V����a��%m�OTz����#:��06�I����n����#"�7�6H@��W��6�ܜE�Oy���Y:�#j�ޟ�Tҟ�JS����`zP��=޹��V�Z��Fe!����ꃇǷ��'Cj�@07�&��#�<C���Y5+\�B���xLs�3�)�=�9��=a�ۜ-;��3�q9�Ќۚ������!s�Ï}���]'=�� �'y�F�m>PZ�!�%�܊n[�˟����Zf�Hږ^�ċ�r=�-P��lbi�5+5e2GǶģE��6���*�U������TDCo��`D� Y!�ܿ�߾S�We�QS��T��0H�qTz��]�U�+�����t[h�e	����3�\���2����u�y�!_�¸n4о�A�VZz��ױ�9�&RsT�G{&e�b�/a����?���q%izy��ի�-�S4&1�Ƨ��H|*���?����O����� F�Tۗ���؄Ą��,]❦���*�ʄg\�2t�a�
>ڍ�2�������$��R-(�I�`�A� A�ԧ \È��	����<j���-��T�l�@�q�ǵ�> 4
���_��
)mfp����Ū .�ߋBI����D`ӯ�`�2��B��2}�o�3Q۲���X �TBT'�i�N�J�_T�`G͹qg��n���,p�x�fs���Y�k˝q�:�N���T��.����j ��to�B�I#RZ�� _�-���������,�7,"';�-����b#ε뺋����f�y���]6T!E�]�tEA'Ż��J;1e��U�4��~�۵�b,H��Ee����E�>�y*w��Ɇ}����������Y2 E��f�5A�b�4�?QqY�gV�c���v��T�J�t����0n�P���q	s{p;5JYB���2>�&5Ϟ��-���	�A�y|�"<��g�m�.[���5���_�̺�2�R*�D��<gr��	�/d��"}�m���9#�$�+�<�?�����k�be����4����Qy�)�a�a������;���u��8��?3X͐��r�����8�E��'D��&A$�[�,?��](������)0�_��h�#�Q���P�Abl����}��ʞ����-ؼ�#d�w�,)Q�wjH�%�1ݫO��@�f��-��tUF:)p����qѬẖ(͒T���,( ���k�n]����O����`؄�D�3�Ғ��P�2����7��_�|<<e[�n���Ih��=e"�$���`�0i����b=ׁ|�m[�/�6�������Q@�4�TYԢy�U-�w-��b~���	�;v��<�W�i�h8�+e�3�@F�V�0��
�R����t-�ݫ��D�,���t�1���)wR_Svx7�T4�����2CK0<���%�9$7�Ք�������➛�k*X1�;��t�L�sg�K18h�Hwma,ߟ,(xH+b�[+�!7�U��|I�T�U6��
ua��v�1O4��O��%v��I=9x[����d�p��z��*��c�ܝu�����^��P�0�s���"�>"�s�V�\�ې2g��ʩ2�_���F 8m�w 5v�1�X����M��X�O�m��f�NgѨ�k�%���w�p�UJ���C�dOCv8y����Zd���[qC�I!�����z�qkYw�n��䜭���<���]	v�G�ڥ��<��]�~{�4�F/o߷���gR'��-��z�i⅟�k��P�`w��?�c E`�!w�ng���[X�ڌ<�k�sP����{)�DAW&尿&��ap��]|!���QǢ\�k���F�T{�6�y��4���|�iCKV����'z(�������~9�wvP4} ��xm��{�&~ Є�p�E~�1j�I+\�7&��	����ry��C$v`hF2b�'y�h\f�n�|�R���#���55~L�}2�nY�����[�_���P������~�m�J�𳜏Zmq`����T��/�
@���[0�s�A�7�%�6}`R��LqiB1� �g��v[�dU�ԩ�i���,J��P<u�1"�|ښb��D��8��\���صtr濧�9�rY��Tg��B&�	���_��i��-�W38���1�k?�5�*��	>��޷��Wd��G���z=���|���������HR�>����+C�?2���8�r�pj�J|ɲ�n�G *p�M� ��w�v���/}b�t�4-L^��#����4� ���0���-�a._�k�Y����$�8������+w�fF�K��£-4��=7��g6<��;�U ^4�������+Z��i�c��5� tb�%��#ACv�!�KҞ��D���i!�����
AiR����9�{wu�X��n'1���!�9)�(����d���H��m$ S�|����i�o�U��[�ѭ}~h�c��Hַ�I�"1�*V_ek��rH#��ü#�_L#�f�SC��&>���'lcKO ���Э�����%�c������?dl�����1��������)��p�����2�w}���As�Xr�����V���}�:��uƕ��w �eX�!s �k�$������G���l�H�
�p�L�'a��X��S��ǜ��8�Wz��|hvz�!�bm6(�4�,�T���{�ܭ�� ��}✃�I�I
{�����2���:;����ZcR��Mo̿�ݞ�p1����f��;�o���9����gS�þl�{Y	=�����<��2��}���)�?�l����,8Z����L����0`��~b���|��8��2>�2���`)Z6m��K��4��ϟS�k:_�~��	G���#��|�t��&��i���k�^5���;*i��(�&X���*�Lk�M��l��5�OU�[}n���|��7�FF'Z��% S��I���ơ��/C"acX������3MVM"ʥ��I�I�u�i�C��
���e��0��{iZn_w帰� �U��ܒ�t^Wu� :����k�Qݒu/چ��m��+����ȜJ;9{�_��@y�\X�۩;/�b���hJ���p=L�_r�(:83n���\th�B�YL�>z� "э�tj�9y��D�/e��� ~�P� L���k|��Es�9|}$�������x�Ͻ{OM����^�au:_�����@}�C}8��K:��t!e �u����6GЏg�G��:�f~��K���4x�u"H-c�f��m��ύ16�I��}&P��tR?F�M�u6��.K�����?���˵�&��bg�b�]<B�q�;�M�J�-������Hۡ}���L��Q��Ц�XO7I���g��� �����0�>_��d���,N8	Uؕy�g
�$N Gn��(~��{�I��!��,`�.Ii�7�W˶����Y	D_�ʼHm��ş����x�f(��5�Dl���0�R{ ��w����ZLY�d��R��q�#ȎJ�r�����0���|@N½.�g���� [q�g����Y+��䜭KF�l����/`����̃��;�(>;����^�w#��΄���{��ʲ����L)�޶�k<̊Ϡ�����w�h�u0 ��,��`О�T�,�=�r�\�MYȧ�&�#�CG�brǒt_���˧U�ofKK���;��Aܐ��"�ImV��Հ���KØ'4s��������ʹQ�xZ'�L=��t�UZ�a���-��ϑ�����Y�,�	VEM�]��k��_��˶���cpQ��@��9���>[̱@im`�b��¬��Z��w�κ8�~�V�aFB�<��U���P�?�&����b}/�Z6ּ����������ml��偹%3J~�(jL:�U����(Cih���x��8��[�a$�1�KB ����KL�u��2���)���4�u�Lݒ��Vh�����2l���ދ�&#�}����P���J�ƶ1��<�X��@�L���w����^��SJ���Y��@�8� ����J��ș��R������Β�k���,���}z�l�_X�W�7�޷J��a�IƬo��R`� �R��ޮ��4�u�o������8_�Fv��B��6���#g͞K	+�v���ό�V'�XA�9�c�?b&&O��s�	`I�wm�R����4x�9X�b���Ǖ��B�ԣPXVƤ�=�h�!�6Z�O��u_�:�����rS��� A��hȍi��[���2s�>��*L��G��sp�Hua�zz�~��2�W�]
~E�f�	4U����������Rh�	¹i��-��t/�����41�lQ�K_dy����1�0��7���=Rc� u���3��z�?�����7�p/�Z���N}Y^����d�]���݆B<I9K�[���q��?�����߉�[�9��>��8ox���D=u)���Q��]j�WT���86��E�<f�����j��7}]�cKk��� _"7�%��gp6LD�*|5)�����~��,gy�8�@���h���;�Y)��"�z`#��㙌VD,t�:@�A �8��-�TԵ�EG ��*J���y���2��^�*c�����}���g�"D=���H�/�z�r$������,�3����	����6(�U�/'t����ި�rۖQ�����z�'�4��D�3GMwT� E:�q�?�'r�e�$�&�ъ1�:X΂V����6$�t�>��`pc�j8 х7x�Ҳ���S|�4�������6�����U��$2��/e�OD+"�o`\��i���*�U��ͺ��~�h��7oP�P�����[�.'y��iS/,g�R;���#����:�,(a�U��u��̥x�#vbٶ@+X7?[��龗�C"�E��,�����1b9����W;^so&'Ft�~�y:���ι�>>=/�V:��Ӝ�P�������	���V�&�	 (-�F'��ph�\f�;)"��R�gH��h(<�z|p�ሳ�Y���թRMl�'�����^N��| �	<���g�Y���?�
k� ����Z�Q֨���=�S�gdd�
g�d�>�ٝ�>��4w�	O9{���C�y���Y��
p��'�`�f￠�%�W�z�t)�@�r�5\{S;�Ϻg2?����u����Ԭ>'��<K�9 g;!��ޒ?������I��������1F�r�|,�0��W�ɯT�{ZgDl��h�x�����s�+�\N�eto��da({����$9�g������]�{AD�?��� �g�aV�,kwH�?�J�� EH']b&��g'��ણX<�`��yD�HB�a�b�>*
��v��Qs̖ؕ�j?�b���ʄ���tڥj�,�\ $j��c�ʛy�rj������p�V��tx�$��|����eޔ���c�bEN�#�F�:��|�ex�L���1�O�r`�EX�9�J�
��u���a�t6��Pa8�%ą�`�;���⻃6kaH#!|�6��F�C�
s�R�F+�E�I�:��Q#������_�I�Mu 	�&��������9KF޻������Uo$I�u�qً��� =e����5��\�Fت�?�4���X�U�r�V�g�X�:���>'f�n0��lvcm G�� Q��g��8�Q�U1?�d���NK*l`\�crn5C
L� 2�ܲ�F�si�{⤧�;����dU���a:���}hc}�|�`���k�/~vϕ���%߰q����Q��������n��u�2�h=q֠�;�Sk.���^Q]%���/���{����m[8*�f�~r)���a���&�~�s��ޠ\vRz���~�2�*�L��,�d{iJp��a���������av2�_dhè4WLf=�n�5׼�ķ��ej:���LoXQP`8J��PO�/|A�>�G{A�P�%����pn�]Y���T��>�����J�_n:������g�����%wWԪ 2]�Ȏ���	a�S���g�|n��ydCXO��Y_�tU<^�u���·&���qd��  �X�K� 2�;ɋ�A�IO�v�0~���Y�����ی�$S�����+�z���Ac��E���s¿cj��j���+��@G�I�c��_��$��0��c��kg��v�b?/�|?��1,.3˧�z��-�n�h���k+�g��h�?��������E�,��������s{|�K��vf8��m�� slE}�Ԥ*�I<�î��y�+��8��r�]�����
p�y��h�숀�Ro�<HYқ��5F����k�Lȴ�B�+�]:�|�����]�S��C13��?���!z}��K�돏~�D��M�Cs<|�'A�}{8_b�!)pB���_?�r��@���6w�>UnS*�?����l����A	8R�*����� ��;B
�k�"���HV�$I\��}��?V�$Y�r ���K�i�P�"�$s�Ia�=�u�e2d���M�y�CI�Q�;C��?8����OK������Ƚ�Xr���B�x��k���փ7o�zM:���^���kZ�E�D���J��py��0<�����jԆWU�� k�n�{�
@J˥6�0ߚ�dވ�&�I2�S@��By}��obtY�B:�\�l�
V'8��
2��_<�PɄ��=$I�����E�ϝRm�aטw��.���rq02-����FQl��A��O�=ꎮ����w���a`О��9��L�P���,�;Gv�'\��h���N� Ǒ���JO��c��j��i�P����d�ozo���������j�a�tF�P,8T҄��CZ��"#BE>�!N�;�)�5�r���j��^ �E~�H�[P�b֒���t%|<a��K'U����9j�.�p�q��"�0F�,G�$]�C�CE��j"=L8�|�y�y.��ly��q�\ho7qא
&6DktAʬp��>g`����4����#��('�hÁ���
&�C%l�=����> #�0�eH����z��
BZ���$m��ƶR2�k��J����m�"���bH��d(3�r�v�\
AP<ǝ�܄�q��`��	|���?W�+n�Ĕ\9���H�Q���Z#u��"�x0�Wė�1d�7OY��*���*pY[��!�0�M�s�}A�Gt���γ� d�7(V��+�9>0=�=4�e*�M��&�{&,��:1
��!�T �Q�8B"��hH���D�"���LΈ幁1R-��ju�rO+cO,6�l�R?\�s�A\h�Z�aD��ˏ���GP[��%�4+CA�Ht��&OpOo�W�,��}����=?h���D �&c^�޴�(�Vrs~��OF�^����0*�}*���4}荶�AI�I|q�S���j�a0AV���^e=n@ 
)г���Gu���'���yK��8�ю���K ��u��-#�	֝ �S��	f4A]/]N�6E\�XZ�Ge��<w#V3�a�	��JI�^$������Жg�]����d���^�RB/�����ta8X�l/��7�-�U��ыKL���G"A4�FJ$I�_Q6�i�y�z��:�K30���:�x�m�,'�ٿ4�e��gV�S��i�	��x��0����B<c@i�Q��4c� 崪}�ñ��\�I��#W��'d��b��	C�������5J:�t�d����G6lʁˏ�>�$%z=�B=�A��G��-�у�Ȣ��_��.��$%�j����Q�I?M&�ϾzB�E�i�tx^��vb'SS6��n>�
����[����n.���D��:��`r����l�$z��Af*�%��w��D����r$|�R|+�vLn{�������.ե�2�~�vɲudfN�9
F���l�x���a�P�E�$�aB���*�E���L�}�8�'h���,[���@Ǚ^�7���t�2"����I�ȉ�ȫN�x���U3Չ��FQ�Q3��0�V�נ�YM�>%O�\��O�"��dl�y�G���z�NR}����f�F���o��;N�aݑ�[,�F�lU�\��k�ѹ,ю��!�D[=3��לx�#��=Y�2�5��`r�5W �Y���E&)~�aN���0"O7`�5+>"tLޖq�Ug�,�gV*[�&h��π�.���Y>����+������g�QL&�n��s���pH]�Mn����jʶ���L��$�[��	�����~�����F�9�ygC-IN��ilc�A����Ϳ�*�&��O_�}#D&�\J9ݩ�"r�Ao@���Qh��Q0���)f���a�f����$|�sfuj��[ÝW��$W�z��k���d�/�������P��������J�G�gŬ���*ݡ�O�v�-�ґh�v,u[���x%��>�6&���|$}@֗��%Gd�49)�ᬒ��s��z��@�r��e���(uI^p�|�T0Ҋ�#	=;鼸�r!�S���N��(4G�����r��=0��V�}�����8%�r��)�nz�x�E��ר���_�7Jq&�on�@"8�D��"�<�y'���B�f���=� !2y��~3�hٖ��i����"���+�ǎN1��!b:T�ne��ǢX�}�4�3���5s>M�$�A��o��c���i�g�e�B2Z)9N����I?U��m��<�����3��rp�5�<��3���`�Y[�c�>=܈�&yOtFpK���r�ܠGH��������)�#���e^�Bѷ(�h�b��؍8R���a�x�V�e��E�	��+�h8|��ɠ��n��Z��S�7�i�LW)��0�,�-{5���� �.�8�,�C,v��,���KuE������3����	����d����?��!���J�l�G'���C�$Z?u5*��p�Z��[��Nװv{ir�7s[\���B��B�z*�p~��	�Qb�6U��� y�T;�ԋ����Ɔ��S�u�����`Y��\�u�w��ŷ��B���5T�Q7������s�F��s��7"���#��|�=M�a^�(�TW��p���3>�n�hk�N'Q�ձ�.P�7��ʟ��l��9]���JGU�c��l�`��+XNA.a������$�k�BO�0*�)r�MB��-)D�}H��[|�:2�3��`IAx�����6���J��Ml<������k��I��і.�t��
���<U2�&qG�6�V�z�1 �����0��|U'Չߔ?����	���̝��^ݽ�&34#D7��cJw���b�ҀW҇��B�V��͙m��}v7�5�>�l:;��N���f=�zeyzG|D�Pu��""���ؚu�3��g��	x|��i�T��s�|X�`cKl�����Tdo|:���A�8['ط�U~�_��:� �y���#�t�#U��C��1�����T- ���=i�J��Φfpb]~���B����z��7l����*�yX�|����"{���<��k�H�W���L����z��\#|�G�8���Y��(�#� &���#�p(X*tY�����3Z8�YFI�T�V�<]�A`}D�U���`b��*J߸�eY��Y��%2N_�4�"�F��s���w���`~I���tx����Xos��&-������
q`Bs8�XX@�P���a��b/�����l�f�{ ��A��r\��`��}��	�[�z�1����߹H����iYk�O�_�D�$j�Iߖ~�+�����lk]n����#�d�6�/�v�E&|Ύ�6�+n���H��QJ��T��b�t?!À�X#
�Be���ޝeW�19/�odq%}�	9U��JL������~ U��'�ʼy<(?a�0�`���a�l��*F�8�c6�~v���*/�׈O⑖���/b�Y�#�,����Vm�=΋��pc��hcx�;M$��NO
��<���ę����#��D�+��l�feԏ�oijZ����S�W��\Qv(� 66\t��Lra��H�y�3�\x)F���]�T�b�ϗ�I���ռ���6���zP��j���SvHeCkrt��%���+\�c11�����(-D���g d��U��I�n�k s	
��Κxϙ撰H!���\�68�%N̛��bkp\"����c����P���� k�4(�nexg]h��r,�>����+8:�a����B��� �,9iS� ��yK�gE�`�O[
`�-C��W��;6�?�A����0N�w���xzoJ�8�].]�lA�hv�Tȍ�PK+)�8O��^�+ �/uP f�{şg���5�U4���M�SgM6����B ��L�y<�9��©Y"���N��$�"��	Wy1΄#&|�f�������c��u����ݩ��[ŷ��A޹puޣɝ������Eu7^?)wy	/�W'h�a�,��^�º>��7 C0�S������1�<�'�B��@^�?u�>���i}�;�u�>&�4"�O�	$�8ZF5a���wx��9�������p�R��s���Xi.S�|��U7m��0����+=9<�{ÁS^�_,��gk�:�LO�	�_E:�ŷ�˳��!�,V�F?��04�Z�N�Ν	Y���U�u�nt�����O��sH0ԫr+;1R�(O4i�\7���t�a!�	�w}��wW|Y���������9�GyL5u��ut�f��q��..�9����&r-1Y��� �~%)�wZ7T���'.a�'�)R���t�ST��r_6tZ�<<Q���f+�2?�c��@D&vG�(�J�P�;���]8P ������u=
<���m�'�I��z�}o�8�[*��&KP����m�� ��n�Ž�������\K���Kzjv��?�$]Qi5���Xs�j�xl5�㸻f�텫�� �^l�O�j �8�B0����zV����Tĵ�}�"����fJ����q�:���ٗ�PAB��R�/	'���/�IlV�+�b������=]27i}�� e�`�Ƕ�D�	��d��s�t]#93�t$<�;�WD�g$��V�]���A���Җ�i�)�*��ꗜ�:�X�oO5��{f�~q�/�Z�i

g4��M�9)8%j�(	(v�_���+�3p"p
y�E��8�����y�Cf[[�=�.ӿ$�ea/ծ�d7wT��v�YN�g�1���~��S JV'd:m�g:��[g2��th[|�I�6��I��z
��Q�'�0P����KN����q����G�p�B�97��	�����"Ԋ����]��V��Z4]�"#��^�U"�Ҍ�3$Z���Ԧ�E^�|uR�)iW�gZjƻY��qP9��W�z��b��-}$.o���������"����$ J��	N���� �����%��tNZz�~�QC��H8XtO\ a��
�-z��u�����_i�cpCz�!Ǔ������g���Y����+�|�������xՅd�x�d�6�ꧧ*�0c�mG�5�/;G;�e����e�pe���f��O���PA��%��WF���|R@wg��@�X�����؀x��Z(X��3$<�x$��S]� ڃ�I&f��h/d�:?��n";?�b��L�y��q��hkd���#�%�Z8n��	����X�]�6�k�#��3y��s'4Պ?r�x����;]�Z���k��8�GT�A��R�H�_�1�I��q�T���환%��Q
����bn�^��7�C{>��R;��bC�@��QQ��Ǿ�x�N:�C�H�Rv-�B�'m>Ӧ�j��#p�R\ΊFk��]��J"ب�I;O��7���z�����-�-�˲���4:b4wS�����!��c{��7ͼ@��Ѐa�p��5Y�dYf���13 ����&������[M��?�Ϲ¬���z!��$6��ċ< �+���v1�˯����ٮ�k�(�3���JJ4��HqV��=//���y�����,��z�]j�m�*2���)(ְ�Yr���Nx��)����&��k���B�����&�����!4�����\����0�ݘcw�	������6a�;�]��~mFh7AIAJ�k���D�"z��C~׾Yy����v��j=ƌ]Q`�^O~d���_`�?�X�K#����ҫʨ�1�R��Vy�NI(�N�t��O��um���f�����pJ�v2���+����g��EH�V�Wz��"��/!J��sD%��7���h���7��b>�W�Oy(���{q�;/�:S�����j�����ia�ۛ�T�6\7m�7!l��t�L�?)x�Jni��;����%&����
�u��3�9tgb�*��N�/b rq�T�>��(�%^Z�������ݴixV�\zX�]����m�d^P!�kb)I����i��l_�f�Y��b�tyntil��By��P�ei��H��a�q�z64_r �F�%C��p7P��c�b]E�Sc	s�D�䩩a?�WX�2���ܸ�ش(2Ë����_J�Շ&(cD�K��cH�Zc �ĺ�P$���F,7?U2�_����@!�A���YiI�"}7���P��#����t7N�@��Xu��E@�����|�ػ�֖��A2{X�_�� ��rUu�B�/��@!Y19QL��� H,�80I(P�o�bЏQ��^�&g���bO/�T/H�q�E�8����a�R#��N���گWN+��B>�&nJ�L�z�?��T������W+��8�����.�P���TP���#D�Vj�\�ԭRB���t{��u1>�	vG�_�=����p�>�gႲZ���X�	�O�8Ԥ�M]F�צ��=~���g݇����� �bE�X��l*���f��a�V�|;���e���;��HBV�_FK]��hI���2���)���Ǖ�a`ҍ����V����3��C�Rt��"� ɼ7�|
T��X��,�A�G�q�ҩc�ũS"�_�I��N�e��Eq�<q[H�S����K�b�"Q�Cs�����Ðm��K1���G�+��?�TCǧT��ɗ �)k�G����,��p��-u�hɖ��:o�%�-c�Y�Q��Ҏ�t��k���ي.,��wӵ����1*�7dO,58��ۜ�Q~��z4R�~��>7�1z@����͚bՖ��H~��N;�Dޯ�J�������K�_w��a�f��d��7b�^"�A��{�({��������C���aC�.�6��r���R!�ՉOA��q��24Q��ϳ[ް�Ĵ�`ZQ��!�"|H2ٟ�?]��-��2�WM���
+���ٹ!�a��ʖ}��25/�Q���,0����0�l��v{9�Ϭ���E���D�؋e!��	�0=�~���ER��~~��w�1E�� C�����=HXˇ������PAmK�k�z%�%����	A�i"h�m��"2$x��y>�R���ϧ&l5N�$�̏n�W�a�Y�M
��fg,{��F�4��3��r�T��!�	Lq�0h8��(�35���-�K�K��ܻ6xD�ee��q$7��[�.��DtL �4�2֨����f4�`	ٚ��SV�ǘ�2�Y�{T����b+�]GyJ�	�
��l;\�2�~o�PWEe�{��Y�P��U���w���S؇]��M ��-�]* ,%�bd 	��ˑd%h�Л�	���6����Y{�2�㿍,�#��qQ��91��d�t9�ۢ�S6��.r�a�g)���oƓ'6�J���*,��T�g�2$�������Jn���L�)�]��2�?��B/U%>w��,^��
�`_k^�-{�l���TV�%�W���S)0����P���Km�G�$���$�Ob��1Gm�e�߃��"�����s#�O^ǈMEQ|�i��̅��\T9��i�����������j�/
{��n�tz��Mrm4�1N��*ndo�����ּ�`|}���j>�� ���c1�ZJe.��{�F�T�6C]pՔ_W#27F�#��]�uTU��D������l-�Ɲ���I$%�?9�G������f&���Q�e�5l�������f�.q�*T
��2�F�ш&,�
�u��u�m��}��z����q�Iq���D�Ѳ��ݝ�9������,r��M�����L�ϵaq\���'M��� ]��{��ubg#�v��-tY�1�i�˧�e7h�i�_��1!�
��KA>��ϙ-�*��⦍0�Q�J�3����\�cxG�����H|ɡ;8e/����r�����n��H-�k�r��@��:����-׉�ミ�ko�f�/��i��pRdz����M�h)����������G+�rgNs�ҟ�Jt�yk�װO�Y!������ּnɅ(�{lP�,gK��cӪ<�;̴n:`L
�m[<�[�q������QS���7�{҃g�����k���mч��o-�? q�W� ��D�|r�A~��2+�bΈ�-���k�����7e���1�{��GU������w6Q��_�+fO
�
�ϑ4�&^��]Y9��5Ht�VzS����B?�-H�s:6_�|�YX����+`1��|nX�[w�bJ�5}��?h��M/�w^�!�^�o�١'�ʒ��2F�1��5����GB9�AO��ǭ��p�Zyc���z9IB�=a:��u��@�WL��g���m��D5Tt�h�q��"�3����ܵR�ʼ0���9EM�>^���g�W�	�d�NIi��#�4��\Uv�O�X�F�xqQ�qH��h�X�C<��]NQ b#Nc�������������(.xQ,�$�M�Z�w�o�(��yS��$��/�q0г��(���Z�%c�I�R��F1�B��;d\��P������Y\Kҝ@��*i�A;7arm��3/í�!�_׵͒��Ɓ�s��D)T\hY�sU��q���*3U�rBZS��v{�Z��ϒ3 o9xlK�\� ?}7���K�� �2�vo����_y�S�	���G�B��z��N�@.��W�����l6��f���ע*\��s
�n�=mXbH�p��&�\�����G��{v@m�\�	}:	t���>��E�r��Bz�(J~(�Q��5�kj�gFK�����f�e� ��G����5l>gX+Y��y�iN��`6.46N\�N�`�Q

�*�p�t���P)�/��������Ȍ�C�Z�D%DD������bf���:9�.dn�Z}U���_�Y�R�o_���R[�V-�Љd0�G�|V`�enekguփ��X��MckV����x��T�:N��/:�#s�8��ǲO(�f����m�EvH����]<*���-;��P�*O���*Fb�j@��ןO鸚����+>�FIsU�����g=��u ����i�㦋�]���hAA`�B1�kC���M���Oy�W��v☔`�%%Nw�Ϻ���L)�g�s�n����	��YRI������}��ie&ꢉ��M�#�VS�e��i��ukQ���XE����jT��1�Q>��mr^좵��}��2��X�zT=��@����ً�Ek����a�]q}��(����]I���y{��3�,+�D5�	v�]����L�x9i-�wy�g��+��^�P�s����֢C ����.��7>�\0E�mfBt �ˠDc�]u�/׬��C~q��d$���l<cFg�����[
S����4�6��5�@��@^��@�^�	�%�z��=���<��rsyw<<k L�&�$iA��lS=?:ˤ�/���+���֣䤯�+�����]�|��g��q*�_�[@(o(�� E[ڤk���J��) R*)b��u���Tk�p5�:��Ы�t$^,v��a��2��_�SsAX�?�,�}n�ӯ{}[�LY������7ƛ�r�m��`&����[�L�')�m��W#���⪟v�P���K�O�Xm�
��bE��:���Wc����C������~��#�UD�s�%�U(�\�Ȗ5�	�5�!�Ɋ}K���Ɔ�R��'g�'7&�O6�
�>��K	�p$�IHԷe��:�a7٪E-��!�l�Y�
��5�P+�����1���giaHǓ�rJ�"ThQe�}^z�1F2݌xz����yu���ߦ���7(�гBo�ok_�M[��n`g�T[��B�G�H��?n����b`)��hRd�?@.b�����M�D�6$��`�	��,R�3ͧ>5%T˪��.���cY=V=xʓ���eW���a��t>�s���j�_�}u^ktA3�k�XY:BK�M�2㢸��y_s���9K� *vFZ�JG��Qyr�Սޝ�Ʊ3۹����5��n�I1�8{�����(�Y�^���|��</�95�=d��a�)%j��
�Ė�,R�I��4�2#���|~.�<� �v��3z�Tz�`Z�]a%L���)��Q���d�Â<bA]�-�Bq�n�e���Y!�|مƜߚ�6
%B �LI�E:��܋�?-yc� �X��81�.�Y�|]����uU9�d,)�p]�M�ٓNh����Y���3���K�0�CziLdĝm�Zɍ���R�w�%3�@T�]?�����U$�)tuP2xA�"��
�;w��S�2��uX�4�ʤe^����:#'��6��I8܀����f�����aL�ɜ�5�s�[��^�C"�YMfW���1�G�kr���!��KM\��8:�7R_2����w5f�|���~�c����=���,�<�~e#K�y����ҡ�/&�U�C�Yz�K��
�ib�{�)�^w�~�g�'g���>$'훑�9o5�q�85l!%�J�aI�'Q�������Re7�X�`���h�D��������׍6�o1Ket@ X�C��!>_�+'����{��Nm��U�R������,sN�������]s�نyF]o�+����o�tM%�f��ven�Qޠ���5���~e��� ���[�?�f�ڹv���7���o�����f"�mN-���!�q�����@�)H"OP� á˫�$�:UX�0`�*���oe{D�����	Բ�i���=�)�ԍ���L3(���M��;����?��R�����|����x_	���£�%W+��aJ�����vH�A�q^� }�e�?o
����!���+L��E�>��J8$ �``�{�ph2��3�@�K�)֬>u�m���=��}Qq��z"��=U��#ٺ./H���>=Cqv5)'~�=��K�$(�b�5ܮ%��3H�pDM�e�<&pw/LnL3NE�<�Ʋ%tQs�� ^�.�O���H���f�����&������,*}?��KU����8�����] �'7�ngak����+�4�G+����a� ����؜8�Ą8x����7�ђ6c����L�F��?��҃�� ��@韖)�j�^�HUcG�	)U�,p��ꯧȉ�w=�����ΤM2�T��y�蝉�U�8	��nR	�Ǔ�0K����X�a��h*q��'&�(wq��.�ܙa�K|��Y���o�)"��<t��(�ޘ��8ƈ����(���F�L7�T�>�Lc�AP���&O���dx��W#/�̇9�s*��!���M��x�� ,�"�A�Ap�����llt1"����`�t�=�F�A!��U�r4����<&1j�d��7ku��u,h�o�h�ҏhS�#��{'w(T�Ҧޮx˜�ӵ�_+T�8.p��zʵ��� �N0I��ֳZ��j��vgb�X\YB{pGB:	��Ε,IG��ƕc�iE�z�D2�S�T�;?����2�-�\��di�hE7�r����v�8�4�X��09<|�Y0�J��5�����__[H"<ŇKW4cak�q�6��z��xF+�K�tc+�[D�p��s�05�?�m�����H��b���?
��b%�b?�E_\5k�醬rayf�`������tL�����	֕����O�;���;�!Z��y�Goy���ˣ,��0��äp��IH�>��^iX��W��\ w�W����k�]%H�oFɏ�ߧ�sD�P��L�3�i��#`�5�F��w��1Z��;(�NyU�'�i��t�M��B�p�`X�*��0v�)e�c�6��K����h�BC̷���|��/X��)���k�;�6J@�(�d����<ޝ2 �Q�&{'P%��f|��v��Xvͥ�m���
��p���I���^�WE׫޷o��60��ӕ�]������\~<����d(����������y���nh��/ّ�Q�t�)1�Vj�>���xV����P6=ު�]�!g�d6jՎ�4$���$�s�8c"K���d�B�P+�''h$.��(�Y�ph,~�����<��z��ʹA�6�\���B�ģ���-z�3�x�Q��k���Ț�ǃm.F!%���*���������]��HZ��F�80[:�p�zP���U_��)8�(P��}R�hF_�z�Ȉa����Ո��l0�:!�6�
�E��t������c1��Z(����X��,vSTH�,�C�X�u=��C�P{�@s�� ��sf�	�=JB���Rw.췕~�Ǯ2]��hT�Mt�&,noO�MI�ܥ�^� �U>��'h���݊<<*y�4Ľ��R5�?Y���L�|��(]`G��.�h�Je�^�$oI�be�)�����K�#�Z�e:�~�S<�(� ��A$�&��*����'����ND�q{'|(���l{s��O���^'��I�i�.��2��ԮRz������D���Oe�^��YQ� ��C�+)�:]��3�E����!p̯C�P�ٹ��j��Frn}���%�<@��Jp%K�l�4j�Y�#w���0�x�(>h��H��B98�4�4�<o{#v�q�x8��(Ҧgk��L`�+P��g<�����|��.���c���;,�A]p����|�T�`�<�^'ER��~�s<�-����7K��gs�����t,ծ/���A��O�AOl(��)�M�֔�7 �p�Z�,�C�5t��e�� v�<��Ĥ�t�Ю�GH0�QIjp������EUf{nIj������:�����E<��HW0�J�< S���L�KgtV���fH�R�"���T8�k�\�u'O�Y���N���J���蟻"���{�e��Y�����`qG�Ѯ��zӳ�݅���x��-��1;rU�\Xj����V�q,��W<~�UD^�f�͘���d}�Z�W�+z%^/��cWMc7�$`�sU��v9RZ��s>ϥfO�;�6�)�,Z$�b���-c�ii�Df�&Œ��̳G���>	�	e�$�����N,�!�^����-R ��Ok��pVN��'!_���o�cs���1B(nr��NW� Lw*<y%�ź���?[�ɕ��I����,���ܹ��F�{!D
1N�pc?u�� |;"l��뭠�p��+�E�M���c̉I�ts�}3_'��>?Cқ4�V��VK�ªħƷ7���-�I�uӯ_9B|c��p(V���)��>̙ &8 �č��+޾P:��3��� |c:�^�U:�KU�چ�i�
������Xo\6��*ꑡ��d��>=�p飋2�[ڃ�@�	g���gS� r�/��~u긑ܾ �Z�f������ɖ$I��v��|T�;)/�E�p��C�}e�r���k���J��ekSu�p�ܶ߉���i1��Bٷb��:�{'��W�E���m4W�`��Ea�����V���\��5��o¡ůk0�����ݽ���,E.�:���,�GO�燔 +l��G~Tϭ�p=�~lΕ�)���ܙ��7Q�6kȄ�͎B	]q��}-��7�1��Y���G9:�W+���d~�����3r�^6���&No=��5z��_�7����0�^5Bq�2�IӍ�ʙx<m,N�z���3��C3i#ǝ�nv���O[�)a�4��q&؋��po�#���̕�� �E%���.��L��R��kj����èЩY,aX���:�([�� gv_s;j�`6$�3u�
��@��a��[�O߼�i����e� %`$�8P��s}����n|�Pi��+�8R7c�Q��8i5S�ƛ�{l�k�M�j�$F���P1�FSf��\�~=g>ʑ?��ӫ|�/�iĚ:��>"4ʩ�l�,�Oo�w%�J�z�ݐe�9�c���O�s��Z
�'w�J���q0�
гfav�/�S8Y�ޱ ��F�����7��v�wg���2Ħ�*�|�ydat05d��l�S�T�m�t�V$��|��İY�p�v8�3D�`����_g��]�����U���^�`�[��]#�a����)��⢄�ô�㽤�`p�
���<$�Q�{�6V��a��Jf�w/RY����� ;x�f�j�^���P�
u���K� ��������t~��p��X�z	��v9�g�����v-�t�>,v�����*�@�1�n�e��6Ɩ��4�#5k��ɸU�I�g �v�f����h��;-k�zƱV�f�����]3ƧW���%�� � ����|Л�����"��>�Sr��p�,6���Jty:@�!�S�𕄓���d�b��F/�fk����.� �&�� Z�x���m��G��iE�E~rԃ0���+�)��~��*ꖧ��;����
bM��f�8�0�������:{�?��l)�V�M3�'s�Kd���p>�����"�lO;��InL��s�6mq�UB *vh���exT��=~����J�=1��4�|fT�q�ဓa���svAf>��y%�:���orir��i�s���1.�KZ��n�����^_G��!�%����X>Y7��d����E3��e����e�x �����������W+H0d�Q�}�jT��~�r=�ы��ӵ��nD�D�h�����6_$�\�L�Ojtʻ�������#�D�^�h��yq��l�t@�+
M�æh��	A�x��i)$
e�����������o����@�qC��taK͐?��UP���9� g\S�+�d:(�*�L$>i؃:&�-K*�0�����ǹ�5�
�r�?:�	����썽�<~ba�r�H �Q��`_��:�nS� aZ���KC��hD9|�Y!��i�г<���ya���[�e��=K�'��2n�kD��N�����.�eoă�p���Gd]�Ro��I$��)�\�o�&"�=�(�Lx�M����d�Z؅G����*��r�=umr���!���j*���h����0�/Мo��>?�����1U0O|�SaMh�X<�,�zj����_z��=�kz���r��)����׉\|Bni����,�<K݉)]�ȳ���4�t&Ǣc�N^�D�M�O�q�x�<%�sI�J��P�Yԭ6�W�յ��-�3�gŇAڼXgA��G\�$�)|������KN��i���q�?�V�A�Y����������r^�Фx���tvW>�^'�2	|�~��;�H֖��F0�0�tF~�j�	���-��&W�A�]��Cf��o�[���穷�ocM�q-WyM�qNc+����6~8P�ϫ����I>?�ZFe�*X�	/��t�V/�ͻ�he�>��;�m)gAi7��M�G����VϬ3̩��&$8���t�6n�-���A)�_�W���UƆo�_"�L�bS��C&���)�;A.���Y��.�oOl��N��2 �,A�|萛E���+�A�E�N=n�2�k� ��?�k
�,po�]��.�V�b��;��K�2HI#¢���SE4P\�%��:VD�B'H*	v����y�F�u��$n��_h����"�����M��G�p��OnX`^�w�jG�"���F��_�aԴ��	<L�V��D=��¢l)�� ��S=�%����V[RѬ<�Dܴ8-3/�����΢���_�?���kLr/<\��)���6��>�$�	8�>���Ԓu3���<�
y�Fb���8����h��~�.d�i�'�ܒ�(x�[�q�[����J�uj����&T��972K-=����
��PB��΁Q1�aZ>3��哒jV���88bS�|/V;������#Z}Oqi�J�8<�0�ǭ��_/�W!��m�������P3)e��&}�*T�{�Z���a�	��!��#�V1��R�o���w�'ֈ<���������ݙ�p?!Se����]�#ƠR{�\��y$<��O�c�`rr07O�%r�VDA6�K#脊x(/���!V?�.�щZ�����B������A��:�Z+rt��*��V�++�Dt��P���YǤ�n��nuj��>�n�k���y g��U_L���)�n#�PaeXDkh��dK5�H�L:�@�w��US�jө���U�!!���惘�'�Ř~��&�ٙ��&u5��%b�[ J�x;׶�83/S���u!��	E^����D`���%�-�R��!=n����p7����lM^}�p����0��v f�S�h�;�S���9R߉������"����k����C�|�0 U�(�i�s���h`ݪN�Ĕ�r�Psz�9����`�=5�������F0A.Z.�h#?�ұW�����EX,UhG�tK,ň��� w~u�iZ����ו��Kf5P�j��!a��m�[�sꮚ ����Vy�ϏN
� O�HU��%xۓ� �ϳ�6�H�T�3�#�4�:	.ܫ/w�Ik�|ی��8�
6׀o�u���L��¼��GB�=�y�����}�x֔4(�����Z���eK�{� Cx\VɐW��@�YQ��?`���F ߻*`�jp�ն,O!�f~��ﳭ�U����5��ʠ�~�jvF>��Y57t���f�:*���Y�yP��&ߦ��~��,�o;��h��.�\�wa��Y�5��"+ �.�ǑX(
q�)}��wl��y�Ni%f�?�5f{�V��я�K��|㪋�!U�����������Z��)Kǰ���(���Px�5�\o<8H�3�d�l�!��Q�v�=��$���ii��Ϙ}�y�f�"4Y�?� ���6Gz��f�6���������4�r��S�F�%�T2��Z�r?Ƭ���8(�8pN��e�PR']���b��^�U8� �~w��2O.hu��w�%Y0w���e]S;���ozz�YI��B��AZ=��uD���^�f�33�X���"W��9�>�%���,�J�_���-������q3� $�_@��O]RV0�g�T#M�p��6���RZN@ �P`KYP��@�h�}iS���:	Q�;@��%�+��&�QR�QM�M��#�U����,����+-�&�@&�QF��E���W%�<�Ry˸��m0�c#��䈒��g|p�qmP��V���L<��clI-%6q���/�ʈ�D3̍4��XC+D$G�o`�y��~�n�q�����L���p6��Ј5�"0/rՊ�i,�~Ϭ�&�L�&|A`6O��.���Z�j/��H C��5G�,�O=ۘoz��W |�tK�sCw���c_��'�l 89?��R� ���C�MѼ���Q�Da�U����B<�fMᨫ-�6����CY�??�-��`�����vl��E���ڇ3.5�E.<�ƎkB����:,��N�h��������	���F$�����?+�f���<-��?i7 \j7��_+Α��ԅ:�n6{�y7]}�� ��`���%%P���h͘�����0��}K0}���L���s�S��z�&�ow/1��UQ��\�{��q���@�g�������Z�,��~��p�[���0oD�oA��:��Ҁ�
�
��MH�8������4ݐ&���-��&����#`���T��~c������Rڬ�"��*��Ogz�Ho�r�*V�#X{h�.X�nc��3<f49�C�7$K^�Az�a��%���5!W�4�i�2v��!�M��Jl�g�^Ք�?�@͑�D�����{�x�~C�=�Us�As�{�z�Y�,�*�ղ��m neO"xΕ;�#�b5���O%�g����#|�k���7�t���ͽpK]��@�<����_a����7����8=����m֘�1���[I�D3�&(v��}��i�{r�w��+(�E�ċB��W �Z�Rs�D��,�2M��67M0��>�g�k�:!Q��g%s�{�&PZ��Y��h8���<���
�o�	��X��	���O�1�'�u�A�U��#���_A2it�2;��KZ��J���n�,���q��?0_2�6]���#v=��s������O����'(CefS�J�9������ӊ�J�u��H<>�l��0��c�LL�'."C:Y�}E�	�;���3x�d�V��9i�!���$��@c���J��W3���J�'�GB�o��j�H��V�������6����L؇r����s8>$aa����eH?,�:�~�����
MP
�F$5�4�+Y j4�\���@�H0KΨ�@6s�WlUn�����y�F�B�*過U��5h�*h�Q��V1�V�5O��ن�|��JgH1c*���sz�J�2����X��u��.w�Û\ն���N����?'庉�יb��8�e�J��w����+�� k�:�Y�����*?0J<Pg�"�����(�!�΁ϰ��)�:c�#է�V,cwj��h��j:�/����\B��˩wH�U'X/Ƶ�P�8��J��0���q�˓��)��H�F�a�T�٩74�w,!�욫�Js��n�� iv�=��"��x�e������u?�eK:����U����)���D/JА�ܠ�(��o;%�ϧ(���U�z���Еf��!	*�>f�����S��6��c5���g��O������!������ηML6�1(���ŷ(�8h�q�a���B��ێ��ˁ��9$�8W(�8tb�.�l���Z�v�W�� x?�l;�6K�J�4E'�P�e���i�%N%0~��4��D�ɠ��&�'��7� wAp�P�^��:�����@����y7r��V�3k��M�z�;T�����#E ��(x0X�
qxh�tw�@ܥ����[W���Y7o���N��0&��y��ݧE���AR�^jE�������}}���i6�Y9L�n{M�pwRV�-+��7��F'^��ϫ!?1ΓU>����sܖ6���H#���>�ȆA#dؘ��*�,,C��恸�ê$8�NC�Wd#�׏=L5�
�����b��|�a��.k,i��$�u��m�c�B��'�w�Dd��?ECF:�#lf���M�,��a'A��ihT֯$�v�y�b��3I���o �8�����h�l9h W�>�5��+��|m`�s[.�t�|h�pD点~J�(mZ���6��(5�qʊ�X�qy"���7�	V\�h�ӟ�8�5O��V`�����Ę���(&PYޘҬ�Z� �@þ^��[#k�EF��!j_�\�?���9���y�d��<���}t���2�(����Y3#�(�1W8�$��O�z����A�M���	IO�HR���2��o�����Zl��HO��|��LH�]�)�����C�� _�[cQiDf;X̂L��)+��<s��eN� ��ɏ��g�&a#+��.Ꭴk4~6���I�G���#	Ep�3x�ƌ��6�r��X�8ioۖ�񱆂[�ݏ�>Z�Y|W���n�J��1�(Q�)H��O7�D�:1��&Uld�Ι�-��bb�׼_���o�oLRA��һ�3�h�?�=�V�T�ф��|���A�X�%�X��j��(�U��i�@�N������0]˗�uI�o��}�E�>�i/�����<�^��*��I�塡���1�����o��>����|o���z�T��IW�fԔ���,-	��\�%��ј'�����C�7�ַ�p(O���ފ��:�U;�ރ�"�ۃa�`1h�ȋ���ϐ`V��x���c��6O�4������� �TL{ �R��b[	R�3�?̠��I$_��%�i~
�@oĥY�9��_�`ۍ�pݰ�/�AS��xn�fB
�آ��W��^��q'+�5�6s��B���"i���-?�u"[���K�/����X�s���Z�A�|�4�yЋ2�W�A�m�p�7\w���J��m�`U������n?-ӸT��	�2��^�sM{u
����&|���� ��?���6�wD��Az�-�f��Mv�UP�V֖��Iho`�{�~fB�QQW�'7s��6��-N����7��S�p����(��ǒnm-�٢s3�@N����+�.�&m&��0!�<UP�G��n�yN!�_��ۥ8�Y��TRb ��2�R�]�F����YD�nDGB�A{�G�&�am�#� �:�``���<ɡe,��T�i"�)X3�ׂx~8�c:Q��C$���ǘ�N
���u͔y�{�9j�I�utX�s�Ñ1�c�xm|�'�,X�;���<Q9�,<��߸�#�}�ժ�؞'��Y�6ym�u�=�va���<�,�[Ǚ�>����4ek������\f.���|�#���������鰠ҷ�3ժo#���W�1lfo�C�WSU(�u$įS���+H�x���mX�܉�16��gmº�Wng�m:l�Y�W���0v��,�iE��F;F��l��pP�å/N�����u�_Q{�!�2��qR3b
��i��f!�W��gks,�W(Լ�cêE���l<���h�i�[���X8Pv�W�l2C��ȵ���22��گaK�_����|��A/����jB�H7$L���zV�tPrd��C�m�^��К�E��T���'�:��SG�/�}�]�����*��`�N��\��A�oJ2��W�xg�-��A-�m&��N��e�3 X}���-�����c��YyE�-�xԧ}��m��t$�=L3��T4W�7塠��1�o`q\рN����p�\�+- qd�7�}����:�;1V��%����mMB[bG@�;D���ԋ�6�� *t��vU���s#G��g�CR�!}����#T��l�MxD��6�X?ӝיI��	�.����H�� �Ep����(��~@Ȳ��5� zcH�����!��'�Ng�I1x��,r��O��>048��9���:�a�n�@L�L�~��r�)�26��`�b9~@<C���7
aGǵ�Hd;�F��)��&���z�5>j�mY�1����q����)V���/�5z�@ѵu{(��#W���N6L���c�hB�Ӑ�;��5� ɒ�s+ޔq�5�>~��r�_�)��'{�'����+��i�҄;&��TE�\8�$ƎH	�c����pK���\�^Y_~1�n	]��֌�Iݔ�n�x;|UW<�Cvm;��у�9�u��=vPCR-�Aq��0YoX)�pafP�����n{������'�%���r��0��-zP K���g*�}"�Ńpe+�0d�Ϊ�y�]���1 �Ody��><=�\�gU&�M�5sT��wQ�����z��\�m|�ׇ���'�}7u}s��/��u��[N����,;��#�SŅ3����FP:3�����U��y=Z� � ��:ۊ�i#8-��SW�	���k�1�gA)���}1��K����6�*�\��^��D"O�z��E��*�׫yƘ'v�0]�d�0�X��KV Ŭ)�����p�W��lϾ�l

4�Б���A'G�K�8�u�H!7�?;�ل�ʴ6���P�e9((�x��\�X�t�,0�[+&�J[��ㄓ���m��d�Lm�#D�V���YՕ!S�.��׬�lX�8}La��NR���t�!���W(��!�d�R >?:k�[t@1�|��r�E�i��Ԧ�����h�	�����<���e��뜒���!
�1#��o󁱝�Y���h�Rq�\/ő��W�=��W�}�vT�k�E�v�N����Q�����'T�^�nI������bb����r�Ŵ�4dRN�-N����moWQ���=��jޤi�dYuu9�$f�QL���6�+Z�^�ϊ���`������r��"2m�bE��m�<� w'wQ�F�T����g٩ l�^��Ƙ���a<F���� zW������&{	~ �v�Cۙ~mY�Ќ��V(Ȭ}�5�qu��45$���u�.wô��!��G�P��$�
ꝡg�5�ݒo�k�[+��#\`�w<�5��<��׏t���
�|�۷x�8�=���9_M���(������P��d��i�$+?�>zT��)n�1��0����c��s��W���eI�W.���Nb����@s�2$��O&"`�p���R:��U���A�9�}��p<���q��~}Q�����6b��r-Q��`9e���0��7Hs�����jա*��D� �+���ྒ�=��%
�\+s�*- k(�-@����qD������%JD��F�y�]��"�<�s�ݗR��������yV��?V�����7(_ҽ�쾧�Jͯ]w�~&Y^���O�n��+
��AQ��q��k)ȎW�I�w��ð����u��C���`�;?ҫ�ƓA��B*@̮Iuc^QE��b���5:V����`i{W�/�	�o�_p����k md3H��^��N���*�0��so�n3�����Q�pC�h�dRt�bz E�Hg�zWFjؙDo��c�ͤ7��-��2rǻf;O�t�n��B~zN��
�S�7n{�1O	7j����#��L�����VO���6�U�g0S��̆�qq˦�d{)?�Q'*���Áy7�k�н<��Ss�����Z��{o/�V�K6LelR�Pw��/0�b"I�R<7s�iݿAߦuN��O�wS�T� k���К���`�􍸉���.��q9p�i�;?�es޿���<6sdNX_���S��/�!:�f^��I� =�t�����g[;������SꆈW����%(JÌ�a����U��!nD���m�)����P�'>~�y �.�i�xM�R��ם5!���02��Q&W	lSC�Y�4�E�?�jE6N�V$��Q-�5%WR��gRo��O��o5Xq[�2�{��N��Wiմ�Ijm*��.��'ͩ�e��*�S�M
�y/BЕ�"\�D6���H��E.�=�z$�k���<�}/�r���:U_E���J|O�S��Ǡ�0-gx�!�9)�l�o�Ѭ��� �� F����.pC�cɍ�`8����1�N�����$ʨ|�3n�I5qg�N����-����t�xY�le$E�[e.$�/�\�w�9p���ӭĈ�rBI���:\���⎭�e^
[5���!	1���_�af`Ѥ%� ,�j��^�
P���(p�'2B��n��?�=L[mZ���¾���нߴ�/�I_� �>_� �0Rv�0+v'�
�S=tF�\�ɺ��9���A�ES94~������C�o�,�-�� ��ʵ,� ?0���� }/�y�'֭��Vj�R��:�j���#
_�V�ٮ�"�%ge�$N ��M��bTc-�&���W�UC����F�O�
iW���31�=V�_�9�YU�y�?(����"t�Y�nxI��y���JleQB*�Z�<���gM�,���!�����v�iTZ���dڕ+��H7-��N5{��N���Ds.ԓ7�I&pZ��F��]�S�ޓ���z4��k],�
:C͘�mT%�`i�ND	ٹy�7����¶�yg|Ki��ٶf���/!m#<��i"���>���E	�7���G�g��[%B*��B,o
�ko�۳�E����R���ϕ�����VM�}��n+��OcS�u�����XB2<�]��f����]n��hǡ��lO]���t׾�6�ۼ1�PdY(3���%���?��!��y �?ۆ�"ol;�ڦE!/�"��i�R�렢$��2n�T	J�"w�~C"m��;��9fa�wQh��w�iF�����u����D^>���^&����_��(���x,`�:Ĺ?��M�P�U����U�^h�	ˍ�px�	uՔȼ&�;�&���H�jb�2#�rs�k0+u
�����՗U�訾�cs��5/.IH�$�A�을�؟��8��F5�����m.�[[�������Xف6;F��Mt���h�Qq�?7
��SM��r=�w���r���"n0M�p;���ݾ�K�ZĂ��n���*����w��x5��qӓq5
��KȲ,xS8t�53&Y9-������.z[��]м�:O��ywML(϶��a�hi71��SJ��[9.�f����$G��y������s�K<�E����UpuiU{)�з�{��9lE�RC ۵^�9��}��A��OV�1SmB<Un��wq(�w��h�}�8]��@iaJSx(����z�=2�cq�TH�9��������/Ep�J�7;1|ե��I��-r£���"�ZU?�$��w&qP�%׭LP&�,����fSɫ[����5��#�r�dz�^����1�t��:|BB��A�{}t�V��(��s��-�l��D�r�g�F�R!���V� �]y`P�����%����=��C,N�ȰX�'�*�y�Do�m��шy�M�YF)N�7��~��T�o�B�6��'X7����TfX�ۀ�Yw�!./��#��1w:��5�1�h�A�[eۭ\��L��81c��ِ�D���\b�����U����鞱���N��)�%o��?����EL�*�UD��  7�x��9Yv!��3�Kw��|`�u���Q��0��[C��_�3�����d�PX4Gݫ2��Ez�M����w7��wLw�	�'��~yL�_������1��WZDN��=4.ƍk��pKCVB����8T�88*�Z��~������~�u�(�=��ާ���[��֔�e��=�
�w���k������D��W��m�W�0�fJ��d`��`r�:Ifb��	���F>�{���&�[j�CY����Ta�_����+s+�d�ib�0��C��߽Y���j!@����j0��V���"dE�dн�����60��+��3�DDȝ�*�?�1�B>X��K��a�a^Aſb5cވ��)�{�{������1��'�����?�`��t>ة�����=��}���.���4��
ICd��6�M���F�p����
�0S��M�W�몆*��G��s3v��Ɗ��)At;�&C�LxY��n6T��5��2�ܭ`e�d�O$ߩX%:?�3��cL����o�����q������p���<U�/�'�ϥ�[n�j����x(9�����!8���
�H��$�ո��Orę��X��`���g|����0	�#>JX���ݿz�k���h�� �Ewz����-�x��F[�N
���ޕS�[���<�1�����9%�B���5&W������'g5@/�@\H3F�ov�3�S�Ǎ=AX�g{~o��T5;�׸nbU㰮�<`�%�I���>������LF����h
5ޑ��}E���L��=�����m�ڃ�w�q��j�����"JՋ4��#- ����x
�d�T�y�I/�D�!�1������t>��a	��l�������pu�i*�c��°P��?�,Q���m��|��d���I��^�r�����b����Ŏ�6@�����D��XHΓ5��'�����m����D]��RQȕe��w��%/X$�j��}�^�u���Ə~�7mKXY�	c���PA�(�%'��b�$��I�źP�551��n6�.�p��У]�I��/��=���ә�!���F~{��.8����ZMD�#:k�-�4�M�cd�p��/j^N��EmyJ�눍b�h�;W%h��K[#f�./�X�u��q�1{ATǻ�0����iߎP�����	�|.D�����z��(I?֏e�[�3�})��|�a�{�Y��Ts�j���Wr�
�� miڨ��cR���� ���G�1� w�}��)	#�lF��4��+�qZBۤ7�DD��>q�y�|�w#ː��;�<��`d>q���x�17�3ҾGN�3��A��#����[\CN1�.�Bbw�-���Y;��w��&@�IUf�e�O[4?O~=,�����`��9�2:[f(��3Q1`�KE�7�\4F��-
�؎MO�C�87x���z���2Ny�!qpײ~�p�%0�4��1܌[x�k����(�J�đ1g�t���ݚNu�Cz���[�6x��p�
�����R([����w���䆺�kٛ� ���?s3�o�o�;~E���@u�H��M���ǈ�"��.s��Ҁc�;E%T��ze��PF�x�,Gi����Xl��
��Z&p�<L ��̺i�g<P�}g�ȁ�f�3�']�qY�7ׇ"�o�Ԅ9���҅$[� WcQ�6���H�T�"E��2�N}/XfT��H�:5��/8�X��:sHy#�����ͥ8�o�|�x�mw�,6���γ��RW0Û}�m���j�AXu�����EG?�|Y�t��h�h/����0�P�q�xH�(<O$�
���o�W�0#�5���,!�o/I��:G�_\���T���^�rL�t���M�J�!�T�Qq��#�&��f�&?/i!|��)�5�����b��s`�F�ҋ{�L���w.����*y����O'��"d(:�L>�SV*M����P�$Sp8������E�M����Y���@�-�-����f>#����SLs���`"�-W�#I����h�[iYznÖ��v�JFm���b����^Bo�ك����ves� �Śwm�t�v��$���a��}�}�p�i��5�s��&��
��[�3�a+��|ߕ|���������������v�o����6��@gY�q�G�A��kO��=F�]-�P�Ҵ�f�G��7a��f�/D�W�7����JX�W
�A��FN��("��M��p�}sV��D^�����D� ʫ^��0�˹w��h#���V�Y�f��*R���j"~�J����/7m���3�.7`F�m�J:H���n�x_��i1�-Ӿ����_B�cx~db�r���!�K�J��T�ߪ�qeV��jb���4�Ӆ�J��=٘}�xR Q�G�/�Z|�{o�����y	���/��T7�����������^�/�sj�3sL�HK��:�l�ߋ�	��:�3!v�[P��J\�lS�-�a��9�����{Z�Ԩ&�CJm�
�6�C�	�|"`4�� m1��Cҕ�d8�SIO�XE�{t\chጭ}���dgX��-���Ӆ�d"�X�0��Ĺ�ae@�贐g��Ǔ.8_� ��Z��f¦a�wj�^��)Bn{\I�Z�Z>�����5�T�j�T����mo�AVX,����οlt�ڴ9U�<�Y;߮8���Pp��yD������,���C5�}�I��<��]"��h�s�'f�1+Q
w�Z����COF˥��-��45f�XL�/����<y����۠>�$�Escr�F�E5�I2K8�(��Ҵß�����/�3�N�����;����nb*��ѕ�Z��r�E��!�3n��{~x������s%�}�\��֮�	��id)�5}g㽧��eG*�;��ʟC���d�����L|�wsP��}�|z���|,�n��#��ςE�C�Y�p��F���.��\��&b��.C��D�"u�M���q]EEj���Ո�t[-��P:�U ���k��}s&W�޼�X��i���F�7�9�����A�Y�V�[	�(/?�9��P�TwW�>��)Zf��ٜ����F�%�R�x�w�A��h��K�u-��O ��Ȼ*�u�˲��o=���WV�HRk`�I���8>(�"���? �]�p��v� �H=�?O�6R�Ɓ �
M��c�ڒ��I&SOF ^��qX��O���
����P[��6A��vpP�X���b�kc����XA(����X�h���E�H��M��:Q D-��BҒ�l�9�%�"
�����ƒ��mo����b�`'��3!1s=�#����#������C�ń��G��	�A��y�"�I!�ncy���ɪَk���@��Q[!�&���hH!�/kZ±搘(���P6��2h�! ���$�_x�B�NЋ8���e���$�$I����E����	��_�M���mO��:s�����~H��"��
=:	�v�Aϗ��'���yq�H^� vM"D��	,o&Vm!Y�����NI�7��
bu>{�-��rT᱿����1Q0���&i���؍cYb/!�¢���&J35�f�q�	�p�ذ\����I�����7�W/&�L��E���&*�ʻ��U��
��U̩��)R	m!���k7�rk�U���1 h��Y�yBR�����!����O���
������❞�H�Vyk�5��M�[_.��ǉ&&ѲF�&��2T`w��-�6���C^��3fo,Xc��p|��rfyC�#�p�]q�J�q�$`1Ȧ'T�B�����2M��鱩���b>[�s ��)%b����,XO��;yc�_8�L�]+ּ� <�o��?�W�(�3�C~C�K�T��.v�,� �g��6��-���g����[#��Hl��D�]^M���t���~���VƲ�(�:�N��R[�.XZzv��&�g��-�#�K�Y�c��*Tk�~t�^��l�]!ϊX���U*hn�_�°�̝�6�> ���rC
鎟�Xu��ɏ���xT����y鑎:������,��L��T>�����6�f����&K����[�1R����B_��<>8{جc�1��x5V�Ŧ�}���f)-�r�R� 4�\�f�HS*��{��
K�%(��c��_�U�e��F�����6�����^�b֊��u]�	9}�bG�VZI;m��g�'�#e�42m�zF
���O
	Z\=3�A���lBĦ�Bg<�*&���e�'	��4}42�F�p��Xqq��w��.6��8� �XQ��/��bl�4~�d{�wnB���;��7\ޠn���F����)�l/x�"QD�Y�4+K/|�[v�p�S����!�Om�f�T��{MI��ۨI	RZ��E�7èqo�����E�qw`��]��:��~[���
�D�$)�<
D%�1V&���v-.�벐��W�
�4��J�s�Z��p�]_�ա�ͩ^jN���k�%E�i��x��)���P��xEX�\o���I�Z�\���1�Ӛ���1;[��>n�NG�6��`�;n'��uF�Myޖ.�����DX�xuK�ܛ�'!�)q�~����,+�53?�O����>E�R��r�Y^��/bу6K�����W��]�c��mT�}�l��w�Fx��%V�v ��^"*$�� W  ����q>�WY�྾�Q���+^���d�B�t���; B�����>����Io��,���� �D�G��L�����ק���q�E�ASn\{�)=�3Xhd�.`�#T�� KX����G���E�Cg[7ĝ���ք��BFB8�!7�E�m[�Ӯ�9�%Dv7��-m�4l�V'z ��>�Z+[���)Ir��ke���Ƶ��l��'�D��_�=M|�r�uIE��@/S|���ED�t0{"�46�����n�y�K�s�>�e��,�ɹW�����}6�C<"���du����J��l��%��-\�"v҄q]�j�p��e����cSR/�6�l�ד?�F�l�H��o��<@=����wc�M��3C��,�0>/�W�ot�^60t�i��k�� Z��*��� 
�	��0.��v�7}�'֫zH��Z�D9Ȋ#��·0�� �A�${{�t��\+t��{Qw���nee�(��ݶ�G$W�;��R�^]k|�;S�H�T���}��M��Eb�?u�ޤQ�y^!=�^W>1����~l/�ck�E�)i~�Y?U}��1���!�r'��uGD�#+jDip��XPNI��7LN�^�̃Ј
:��VV�4�H1�cCOT���s��#��}�g!k`H_%E���(L1�k}�2L	��l����O�J����B:�j�����Ŏ^SN��b`_v�4?��0G�O�/�X��A�׆�Dp��E��m��V8�Hq-G=䑹�U�N��<��(.����D�|��D���4ǲzI�6k챡)$��7�0�~YU�'�U%�$�K��O����8{C8�"|��h،�%sTrv,f%ob9CC.����օy��~��j��������S_�TE�d����Ȧ��|�_FK����8��נ_?a+����h��8������GAX�:'��x?�������e��J�Qۻ�~ܐ���H^y�u��Ә�>��/:Aq6����jl�j�#����s�8OX�"��O�y!���e"��c�G��I�$���=3��܅D=v�e	�p0.q���N�WM7��A9*o��8 d�%" ���(� Ȱ	�{�x3ùhy%#�j�Mf��mc�`����Nf5���=��:U-x� �w�c�x����Y���DT��x�����ϟ�֌��,�޹�oqa���TI�ȹ|L��lK������d����$rnm� �r�������;��ƥ
;Uam{���1h���ͽ����蝳�W�Sm��ٱ�l�#LP��9��qoL��;Mא���^�A�j~:ײ��V��؆�X���AV����֜S0GS���H��-u��eE��d4�7�??���kh@T���?���U}q�B�PX�N��/ 8g�k����k����22�d��蕅`�j�+���.<�?7n5��?���.��������^-���/~!3U��E(�9.
%�$��C�8�y�BP�C1y�A�I�&�n^1��o2	Ħ���vD�+��t�|,�6���ZI�����z��W휭x�'R��8W+�tE�Uӭ�6�&��?� -|�Y|� 3YÉ��͖��f�>�F�1�r�x��);tsO������M��pV�������+�g	%`����L�]�ȔkgA+q8E�x_����eՇ$���t���A~�*�ŭ �n"%�k��Z��Kt6�"�����R��~.^+g�rg���N؇�7��H�M1���T{�����'7�89A	�"���->�AĥJ�|��
>�q�}LHVS;t���DS���J�_j�8�b�o����:��Z��h�5��Z�\��
�>p"Ο&�����g�mi���	Q��� AYM��`m��	^�EH���>l� :s�A��Ax#t���؞�k���$�%J�����%:L}����vo�� �w�,Dc}X����ZlaX�"��t�b��t���HϿ��d(i��<�x��G8�ڔ�dG�xڠ�1�M�2�U!��+��!}p�:����� ^;�K�b^�|Y�u�wh��?�i7`���zA��x��ʄ�T���
�V�8#u�цE�6:��uS5��vSe79q%21jS#�^䡠:��?b<�e���p	�$��܆p�g������MSg/;X
�u(6jb��?!��5��{XT�{|Ox
�,��XL��& Pv�a�X�6�7k����n��*0aW�R���NN��s3��q#�f!4�TD��(ntU�
�O���y�疋��4*}Rˆ�fTj}�R��Uk�C�eiv7N�,�8�MJ�M���$n�֢�E�t|tP�� ���x����ő�+��~a7b�p�O`i��#����Ǎ0A���Tg���v��
�6��ʍ$�M���o���������Z�E��a�C0�/���#�%�X?7�Y�|.WMF}�-��@��Z�-���G�<���`M�N�������+V��϶8��e1SBTw͐�$ʻ!�������v���R9%{_��s��D���O��՜m�3n'~j+c?ʁ�z.7��@J��.�8�h�E,1��Z��:���#c�KV���1P��ozcTVL���/"	j�K�}~k�h����P�I�ᒅV��1��F�M�;`�]�]f��S��(�q
 ��ml1QԬ�����hx����4�1�a4����҇��J�?]:z������=u��&N����U5�AbB�+��֋�R�
��te��=�I��������*�U��a㢚�M���Ye�X8�cݱi�!"F��Lח8�׺���;�S�����]k-N�BV|J�F�܄�t4u��DQ�f��$�3J_�)|O[��޿�(�~��{J��c�d���30U�qY��9��>F5�F��sd�r���k�x\G����\�j�}�w �Ye��Q0�@�x*�}�m��5�#�&���ܩe�̉����˛l���a��d�����Ala�"Z��#T���Jb�mI��71��"���p�[j����
 %�T@EƇo�t�I�j�E�&��+��Q뷔�{���f��Ă�)�C�w���iτ*͑����M ���ʹ:����5��C!�{�WX|3Id�?���qwn��˶�,���i-]����]&b�9g�M�Z;���"AḲ�!�$ٮu鎠K����^0� w��E����_O@_Y\Xo�xka)x���$���O���pZ����1�r�ɍ���L����U�)��G�:M� �dXk��ŗ �`��J=�n�E������Bғ��W3t����j�8��?
�d�\͜�T�3�+Ip2�M�m����>������-6%���:�Tӫ[�_���ς�5T|�Sj*���)�3�w�������[y1�ޥ|����;}�BCw*�7G�,#�B��E�&2Xӟ�m�!?����΄z@-˹A[�Fd���UƐ��f	K��[�#��Bz�#�k��d(����Y|#���`26��"fH�߻>ߒ�ȁ3-��2(�-E��Y��8�0��s�L��J@Z|z*���6k���֌�
'�e[�d8
�ϒ��f���� J������X������D��f����|iv���97^T2S���a/Ƃ����'N����6���������
�x�E���	�(�JɜDIvꍽ����;�"ɵ�Mp�@�5����S�������3��L.�1 y:�tB8;����0	��>s7L�:l�̸��4ɟ��%.��8��z�����݇�nk�=�$~Nz�ӊ%��"b��E7J����,���(�� �r �폘v��Lu���G��δ�s ��A7�X����>��ЕU>��fb?��&``��A}pq,�@S���F�2)�Q��w���b�4LgL�UG8v�Q�|!{#h�6%�-��U5��1�5lD����eҐ3P��l8*/��-�	x�7p���U!J�]�0irR����W����48�L��G�o��V�=�I�C:�����^7M|YoӷD����c�+f�Go�?�QK*�ݲ0B�n���Yv[{=h~3!�]�<���ү�◬�*<F�Eh[�?(��?�fXw�p�H3VGӜ��Հ;���wږs�#�7�N�wiT�.��U�[���������cz|.#��F��sS�)�(�����H��w�3�ś*ƈ?�����6��!�� ���3W�/����^�UTv
�1.�����ݔ��X���1aa�;���:���1G.�ꭹ��e�,����}���2��-̈́7Q��%��k�@�g��r��,`��Ͷ&o	�~!��r
#���wY��%^��� x����L_�2q���C�a5�p�/qR��v�_�z���e��^��s�& i�fd5�����Lܼ)��Y�@pDN��˅��q��8%ŀ֔�ǽ�_�N���-��)�2�k96A�~�+~F�%�Ut��Y��]���F"R�k��!Z��}��c���lGC�OϪT=Y���+�$z�I�����sHs�9e}4d��ѹ��NfH�{Zt�� ��%��[�Zb�u�R=kK'�U-�W�+m/d����<	�d�N聛�2�{r��䑢eYN3��[��\ʏz��Z	�Є�rQk(n[��t�p���S�s+�ʸ��G`F6�=>A~� Tp{#�Q}f7Li���;"�Tga�������Љ�{�8Ք	1��|�E����6�_P�I:-w��5��gY�~M�:��&#� ��B���8�vS�6���/�ݝiG0�X��1��}倹�:D����#��剘R?��u[�Hܓ�0�g�ii�:��:������v�b#&�V[�nI�1u�:98��X��z�HL˓�xt����T�����.i�QR��-*"��ZT}�������,4�M�p��T�r3�����1Iq��BEI*9��6s* �Ǐ�Z���rYVWƽH�#% nԉ�Ł��!2�FנƮC�c�I�`�EB���^`�|��0L��`���0M[�hXzgX󜜔�-=��%L���2ާ��#�oAǘ+�U_
 � ;���Y�D���h�W�����cd�3_NK��7o�s#kae@Q���>3%<��_�J���0��A�QwV�i��K؀"*��κb0~�S�V